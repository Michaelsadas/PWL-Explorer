module PE(
  input        clock,
  input  [7:0] io_inR,
  input  [7:0] io_inD,
  output [7:0] io_outL,
  output [7:0] io_outU,
  input        io_dir,
  input        io_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] reg_; // @[Reg.scala 15:16]
  assign io_outL = reg_; // @[Transposer.scala 113:13]
  assign io_outU = reg_; // @[Transposer.scala 112:13]
  always @(posedge clock) begin
    if (io_en) begin // @[Reg.scala 16:19]
      if (~io_dir) begin // @[Transposer.scala 110:28]
        reg_ <= io_inR;
      end else begin
        reg_ <= io_inD;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AlwaysOutTransposer(
  input        clock,
  input        reset,
  output       io_inRow_ready,
  input        io_inRow_valid,
  input  [7:0] io_inRow_bits_0,
  input  [7:0] io_inRow_bits_1,
  input  [7:0] io_inRow_bits_2,
  input  [7:0] io_inRow_bits_3,
  output [7:0] io_outCol_bits_0,
  output [7:0] io_outCol_bits_1,
  output [7:0] io_outCol_bits_2,
  output [7:0] io_outCol_bits_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pes_0_0_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_0_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_0_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_0_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_0_io_outU; // @[Transposer.scala 116:37]
  wire  pes_0_0_io_dir; // @[Transposer.scala 116:37]
  wire  pes_0_0_io_en; // @[Transposer.scala 116:37]
  wire  pes_0_1_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_1_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_1_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_1_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_1_io_outU; // @[Transposer.scala 116:37]
  wire  pes_0_1_io_dir; // @[Transposer.scala 116:37]
  wire  pes_0_1_io_en; // @[Transposer.scala 116:37]
  wire  pes_0_2_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_2_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_2_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_2_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_2_io_outU; // @[Transposer.scala 116:37]
  wire  pes_0_2_io_dir; // @[Transposer.scala 116:37]
  wire  pes_0_2_io_en; // @[Transposer.scala 116:37]
  wire  pes_0_3_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_3_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_3_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_3_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_0_3_io_outU; // @[Transposer.scala 116:37]
  wire  pes_0_3_io_dir; // @[Transposer.scala 116:37]
  wire  pes_0_3_io_en; // @[Transposer.scala 116:37]
  wire  pes_1_0_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_0_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_0_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_0_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_0_io_outU; // @[Transposer.scala 116:37]
  wire  pes_1_0_io_dir; // @[Transposer.scala 116:37]
  wire  pes_1_0_io_en; // @[Transposer.scala 116:37]
  wire  pes_1_1_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_1_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_1_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_1_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_1_io_outU; // @[Transposer.scala 116:37]
  wire  pes_1_1_io_dir; // @[Transposer.scala 116:37]
  wire  pes_1_1_io_en; // @[Transposer.scala 116:37]
  wire  pes_1_2_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_2_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_2_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_2_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_2_io_outU; // @[Transposer.scala 116:37]
  wire  pes_1_2_io_dir; // @[Transposer.scala 116:37]
  wire  pes_1_2_io_en; // @[Transposer.scala 116:37]
  wire  pes_1_3_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_3_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_3_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_3_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_1_3_io_outU; // @[Transposer.scala 116:37]
  wire  pes_1_3_io_dir; // @[Transposer.scala 116:37]
  wire  pes_1_3_io_en; // @[Transposer.scala 116:37]
  wire  pes_2_0_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_0_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_0_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_0_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_0_io_outU; // @[Transposer.scala 116:37]
  wire  pes_2_0_io_dir; // @[Transposer.scala 116:37]
  wire  pes_2_0_io_en; // @[Transposer.scala 116:37]
  wire  pes_2_1_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_1_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_1_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_1_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_1_io_outU; // @[Transposer.scala 116:37]
  wire  pes_2_1_io_dir; // @[Transposer.scala 116:37]
  wire  pes_2_1_io_en; // @[Transposer.scala 116:37]
  wire  pes_2_2_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_2_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_2_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_2_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_2_io_outU; // @[Transposer.scala 116:37]
  wire  pes_2_2_io_dir; // @[Transposer.scala 116:37]
  wire  pes_2_2_io_en; // @[Transposer.scala 116:37]
  wire  pes_2_3_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_3_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_3_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_3_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_2_3_io_outU; // @[Transposer.scala 116:37]
  wire  pes_2_3_io_dir; // @[Transposer.scala 116:37]
  wire  pes_2_3_io_en; // @[Transposer.scala 116:37]
  wire  pes_3_0_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_0_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_0_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_0_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_0_io_outU; // @[Transposer.scala 116:37]
  wire  pes_3_0_io_dir; // @[Transposer.scala 116:37]
  wire  pes_3_0_io_en; // @[Transposer.scala 116:37]
  wire  pes_3_1_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_1_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_1_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_1_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_1_io_outU; // @[Transposer.scala 116:37]
  wire  pes_3_1_io_dir; // @[Transposer.scala 116:37]
  wire  pes_3_1_io_en; // @[Transposer.scala 116:37]
  wire  pes_3_2_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_2_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_2_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_2_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_2_io_outU; // @[Transposer.scala 116:37]
  wire  pes_3_2_io_dir; // @[Transposer.scala 116:37]
  wire  pes_3_2_io_en; // @[Transposer.scala 116:37]
  wire  pes_3_3_clock; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_3_io_inR; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_3_io_inD; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_3_io_outL; // @[Transposer.scala 116:37]
  wire [7:0] pes_3_3_io_outU; // @[Transposer.scala 116:37]
  wire  pes_3_3_io_dir; // @[Transposer.scala 116:37]
  wire  pes_3_3_io_en; // @[Transposer.scala 116:37]
  reg [1:0] counter; // @[Transposer.scala 117:24]
  reg  dir; // @[Transposer.scala 118:20]
  wire  _T = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  wire  _T_16 = ~dir; // @[Transposer.scala 142:29]
  wire [7:0] left_out_0 = pes_0_0_io_outL; // @[Transposer.scala 139:25 Transposer.scala 139:25]
  wire [7:0] up_out_0 = pes_0_0_io_outU; // @[Transposer.scala 140:23 Transposer.scala 140:23]
  wire [7:0] left_out_1 = pes_1_0_io_outL; // @[Transposer.scala 139:25 Transposer.scala 139:25]
  wire [7:0] up_out_1 = pes_0_1_io_outU; // @[Transposer.scala 140:23 Transposer.scala 140:23]
  wire [7:0] left_out_2 = pes_2_0_io_outL; // @[Transposer.scala 139:25 Transposer.scala 139:25]
  wire [7:0] up_out_2 = pes_0_2_io_outU; // @[Transposer.scala 140:23 Transposer.scala 140:23]
  wire [7:0] left_out_3 = pes_3_0_io_outL; // @[Transposer.scala 139:25 Transposer.scala 139:25]
  wire [7:0] up_out_3 = pes_0_3_io_outU; // @[Transposer.scala 140:23 Transposer.scala 140:23]
  wire [1:0] _T_24 = 2'h3 - 2'h1; // @[Util.scala 13:22]
  wire [1:0] _T_26 = _T_24 + 2'h1; // @[Util.scala 13:26]
  wire [1:0] _T_31 = 2'h3 - counter; // @[Util.scala 13:57]
  wire [1:0] _T_33 = 2'h1 - _T_31; // @[Util.scala 13:48]
  wire [1:0] _T_35 = _T_33 - 2'h1; // @[Util.scala 13:62]
  wire [1:0] _T_37 = counter + 2'h1; // @[Util.scala 13:71]
  PE pes_0_0 ( // @[Transposer.scala 116:37]
    .clock(pes_0_0_clock),
    .io_inR(pes_0_0_io_inR),
    .io_inD(pes_0_0_io_inD),
    .io_outL(pes_0_0_io_outL),
    .io_outU(pes_0_0_io_outU),
    .io_dir(pes_0_0_io_dir),
    .io_en(pes_0_0_io_en)
  );
  PE pes_0_1 ( // @[Transposer.scala 116:37]
    .clock(pes_0_1_clock),
    .io_inR(pes_0_1_io_inR),
    .io_inD(pes_0_1_io_inD),
    .io_outL(pes_0_1_io_outL),
    .io_outU(pes_0_1_io_outU),
    .io_dir(pes_0_1_io_dir),
    .io_en(pes_0_1_io_en)
  );
  PE pes_0_2 ( // @[Transposer.scala 116:37]
    .clock(pes_0_2_clock),
    .io_inR(pes_0_2_io_inR),
    .io_inD(pes_0_2_io_inD),
    .io_outL(pes_0_2_io_outL),
    .io_outU(pes_0_2_io_outU),
    .io_dir(pes_0_2_io_dir),
    .io_en(pes_0_2_io_en)
  );
  PE pes_0_3 ( // @[Transposer.scala 116:37]
    .clock(pes_0_3_clock),
    .io_inR(pes_0_3_io_inR),
    .io_inD(pes_0_3_io_inD),
    .io_outL(pes_0_3_io_outL),
    .io_outU(pes_0_3_io_outU),
    .io_dir(pes_0_3_io_dir),
    .io_en(pes_0_3_io_en)
  );
  PE pes_1_0 ( // @[Transposer.scala 116:37]
    .clock(pes_1_0_clock),
    .io_inR(pes_1_0_io_inR),
    .io_inD(pes_1_0_io_inD),
    .io_outL(pes_1_0_io_outL),
    .io_outU(pes_1_0_io_outU),
    .io_dir(pes_1_0_io_dir),
    .io_en(pes_1_0_io_en)
  );
  PE pes_1_1 ( // @[Transposer.scala 116:37]
    .clock(pes_1_1_clock),
    .io_inR(pes_1_1_io_inR),
    .io_inD(pes_1_1_io_inD),
    .io_outL(pes_1_1_io_outL),
    .io_outU(pes_1_1_io_outU),
    .io_dir(pes_1_1_io_dir),
    .io_en(pes_1_1_io_en)
  );
  PE pes_1_2 ( // @[Transposer.scala 116:37]
    .clock(pes_1_2_clock),
    .io_inR(pes_1_2_io_inR),
    .io_inD(pes_1_2_io_inD),
    .io_outL(pes_1_2_io_outL),
    .io_outU(pes_1_2_io_outU),
    .io_dir(pes_1_2_io_dir),
    .io_en(pes_1_2_io_en)
  );
  PE pes_1_3 ( // @[Transposer.scala 116:37]
    .clock(pes_1_3_clock),
    .io_inR(pes_1_3_io_inR),
    .io_inD(pes_1_3_io_inD),
    .io_outL(pes_1_3_io_outL),
    .io_outU(pes_1_3_io_outU),
    .io_dir(pes_1_3_io_dir),
    .io_en(pes_1_3_io_en)
  );
  PE pes_2_0 ( // @[Transposer.scala 116:37]
    .clock(pes_2_0_clock),
    .io_inR(pes_2_0_io_inR),
    .io_inD(pes_2_0_io_inD),
    .io_outL(pes_2_0_io_outL),
    .io_outU(pes_2_0_io_outU),
    .io_dir(pes_2_0_io_dir),
    .io_en(pes_2_0_io_en)
  );
  PE pes_2_1 ( // @[Transposer.scala 116:37]
    .clock(pes_2_1_clock),
    .io_inR(pes_2_1_io_inR),
    .io_inD(pes_2_1_io_inD),
    .io_outL(pes_2_1_io_outL),
    .io_outU(pes_2_1_io_outU),
    .io_dir(pes_2_1_io_dir),
    .io_en(pes_2_1_io_en)
  );
  PE pes_2_2 ( // @[Transposer.scala 116:37]
    .clock(pes_2_2_clock),
    .io_inR(pes_2_2_io_inR),
    .io_inD(pes_2_2_io_inD),
    .io_outL(pes_2_2_io_outL),
    .io_outU(pes_2_2_io_outU),
    .io_dir(pes_2_2_io_dir),
    .io_en(pes_2_2_io_en)
  );
  PE pes_2_3 ( // @[Transposer.scala 116:37]
    .clock(pes_2_3_clock),
    .io_inR(pes_2_3_io_inR),
    .io_inD(pes_2_3_io_inD),
    .io_outL(pes_2_3_io_outL),
    .io_outU(pes_2_3_io_outU),
    .io_dir(pes_2_3_io_dir),
    .io_en(pes_2_3_io_en)
  );
  PE pes_3_0 ( // @[Transposer.scala 116:37]
    .clock(pes_3_0_clock),
    .io_inR(pes_3_0_io_inR),
    .io_inD(pes_3_0_io_inD),
    .io_outL(pes_3_0_io_outL),
    .io_outU(pes_3_0_io_outU),
    .io_dir(pes_3_0_io_dir),
    .io_en(pes_3_0_io_en)
  );
  PE pes_3_1 ( // @[Transposer.scala 116:37]
    .clock(pes_3_1_clock),
    .io_inR(pes_3_1_io_inR),
    .io_inD(pes_3_1_io_inD),
    .io_outL(pes_3_1_io_outL),
    .io_outU(pes_3_1_io_outU),
    .io_dir(pes_3_1_io_dir),
    .io_en(pes_3_1_io_en)
  );
  PE pes_3_2 ( // @[Transposer.scala 116:37]
    .clock(pes_3_2_clock),
    .io_inR(pes_3_2_io_inR),
    .io_inD(pes_3_2_io_inD),
    .io_outL(pes_3_2_io_outL),
    .io_outU(pes_3_2_io_outU),
    .io_dir(pes_3_2_io_dir),
    .io_en(pes_3_2_io_en)
  );
  PE pes_3_3 ( // @[Transposer.scala 116:37]
    .clock(pes_3_3_clock),
    .io_inR(pes_3_3_io_inR),
    .io_inD(pes_3_3_io_inD),
    .io_outL(pes_3_3_io_outL),
    .io_outU(pes_3_3_io_outU),
    .io_dir(pes_3_3_io_dir),
    .io_en(pes_3_3_io_en)
  );
  assign io_inRow_ready = 1'h1; // @[Transposer.scala 137:18]
  assign io_outCol_bits_0 = ~dir ? $signed(left_out_0) : $signed(up_out_0); // @[Transposer.scala 142:24]
  assign io_outCol_bits_1 = ~dir ? $signed(left_out_1) : $signed(up_out_1); // @[Transposer.scala 142:24]
  assign io_outCol_bits_2 = ~dir ? $signed(left_out_2) : $signed(up_out_2); // @[Transposer.scala 142:24]
  assign io_outCol_bits_3 = ~dir ? $signed(left_out_3) : $signed(up_out_3); // @[Transposer.scala 142:24]
  assign pes_0_0_clock = clock;
  assign pes_0_0_io_inR = pes_0_1_io_outL; // @[Transposer.scala 123:26]
  assign pes_0_0_io_inD = pes_1_0_io_outU; // @[Transposer.scala 129:26]
  assign pes_0_0_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_0_0_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_0_1_clock = clock;
  assign pes_0_1_io_inR = pes_0_2_io_outL; // @[Transposer.scala 123:26]
  assign pes_0_1_io_inD = pes_1_1_io_outU; // @[Transposer.scala 129:26]
  assign pes_0_1_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_0_1_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_0_2_clock = clock;
  assign pes_0_2_io_inR = pes_0_3_io_outL; // @[Transposer.scala 123:26]
  assign pes_0_2_io_inD = pes_1_2_io_outU; // @[Transposer.scala 129:26]
  assign pes_0_2_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_0_2_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_0_3_clock = clock;
  assign pes_0_3_io_inR = io_inRow_bits_0; // @[Transposer.scala 123:26]
  assign pes_0_3_io_inD = pes_1_3_io_outU; // @[Transposer.scala 129:26]
  assign pes_0_3_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_0_3_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_1_0_clock = clock;
  assign pes_1_0_io_inR = pes_1_1_io_outL; // @[Transposer.scala 123:26]
  assign pes_1_0_io_inD = pes_2_0_io_outU; // @[Transposer.scala 129:26]
  assign pes_1_0_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_1_0_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_1_1_clock = clock;
  assign pes_1_1_io_inR = pes_1_2_io_outL; // @[Transposer.scala 123:26]
  assign pes_1_1_io_inD = pes_2_1_io_outU; // @[Transposer.scala 129:26]
  assign pes_1_1_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_1_1_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_1_2_clock = clock;
  assign pes_1_2_io_inR = pes_1_3_io_outL; // @[Transposer.scala 123:26]
  assign pes_1_2_io_inD = pes_2_2_io_outU; // @[Transposer.scala 129:26]
  assign pes_1_2_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_1_2_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_1_3_clock = clock;
  assign pes_1_3_io_inR = io_inRow_bits_1; // @[Transposer.scala 123:26]
  assign pes_1_3_io_inD = pes_2_3_io_outU; // @[Transposer.scala 129:26]
  assign pes_1_3_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_1_3_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_2_0_clock = clock;
  assign pes_2_0_io_inR = pes_2_1_io_outL; // @[Transposer.scala 123:26]
  assign pes_2_0_io_inD = pes_3_0_io_outU; // @[Transposer.scala 129:26]
  assign pes_2_0_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_2_0_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_2_1_clock = clock;
  assign pes_2_1_io_inR = pes_2_2_io_outL; // @[Transposer.scala 123:26]
  assign pes_2_1_io_inD = pes_3_1_io_outU; // @[Transposer.scala 129:26]
  assign pes_2_1_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_2_1_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_2_2_clock = clock;
  assign pes_2_2_io_inR = pes_2_3_io_outL; // @[Transposer.scala 123:26]
  assign pes_2_2_io_inD = pes_3_2_io_outU; // @[Transposer.scala 129:26]
  assign pes_2_2_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_2_2_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_2_3_clock = clock;
  assign pes_2_3_io_inR = io_inRow_bits_2; // @[Transposer.scala 123:26]
  assign pes_2_3_io_inD = pes_3_3_io_outU; // @[Transposer.scala 129:26]
  assign pes_2_3_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_2_3_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_3_0_clock = clock;
  assign pes_3_0_io_inR = pes_3_1_io_outL; // @[Transposer.scala 123:26]
  assign pes_3_0_io_inD = io_inRow_bits_0; // @[Transposer.scala 129:26]
  assign pes_3_0_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_3_0_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_3_1_clock = clock;
  assign pes_3_1_io_inR = pes_3_2_io_outL; // @[Transposer.scala 123:26]
  assign pes_3_1_io_inD = io_inRow_bits_1; // @[Transposer.scala 129:26]
  assign pes_3_1_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_3_1_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_3_2_clock = clock;
  assign pes_3_2_io_inR = pes_3_3_io_outL; // @[Transposer.scala 123:26]
  assign pes_3_2_io_inD = io_inRow_bits_2; // @[Transposer.scala 129:26]
  assign pes_3_2_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_3_2_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  assign pes_3_3_clock = clock;
  assign pes_3_3_io_inR = io_inRow_bits_3; // @[Transposer.scala 123:26]
  assign pes_3_3_io_inD = io_inRow_bits_3; // @[Transposer.scala 129:26]
  assign pes_3_3_io_dir = dir; // @[Transposer.scala 133:32]
  assign pes_3_3_io_en = io_inRow_ready & io_inRow_valid; // @[Decoupled.scala 40:37]
  always @(posedge clock) begin
    if (reset) begin // @[Transposer.scala 117:24]
      counter <= 2'h0; // @[Transposer.scala 117:24]
    end else if (_T) begin // @[Transposer.scala 144:24]
      if (counter >= _T_26) begin // @[Util.scala 13:10]
        counter <= _T_35;
      end else begin
        counter <= _T_37;
      end
    end
    if (reset) begin // @[Transposer.scala 118:20]
      dir <= 1'h0; // @[Transposer.scala 118:20]
    end else if (counter == 2'h3 & _T) begin // @[Transposer.scala 148:49]
      dir <= _T_16; // @[Transposer.scala 149:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dir = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_16(
  input        clock,
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  input  [7:0] io_in_d,
  output [7:0] io_out_a,
  output [7:0] io_out_b,
  output [7:0] io_out_c,
  input        io_in_control_dataflow,
  input        io_in_control_propagate,
  input  [3:0] io_in_control_shift,
  output       io_out_control_dataflow,
  output       io_out_control_propagate,
  output [3:0] io_out_control_shift,
  input  [2:0] io_in_id,
  output [2:0] io_out_id,
  input        io_in_last,
  output       io_out_last,
  input        io_in_valid,
  output       io_out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] c1; // @[PE.scala 50:15]
  reg [15:0] c2; // @[PE.scala 51:15]
  reg  last_s; // @[Reg.scala 15:16]
  wire  flip = last_s != io_in_control_propagate; // @[PE.scala 68:21]
  wire [3:0] shift_offset = flip ? io_in_control_shift : 4'h0; // @[PE.scala 69:25]
  wire [15:0] _T_4 = $signed(c1) >>> shift_offset; // @[PE.scala 82:23]
  wire  _T_5 = $signed(_T_4) > 16'sh7f; // @[Arithmetic.scala 126:33]
  wire  _T_6 = $signed(_T_4) < -16'sh80; // @[Arithmetic.scala 126:60]
  wire [15:0] _T_7 = _T_6 ? $signed(-16'sh80) : $signed(_T_4); // @[Mux.scala 98:16]
  wire [15:0] _T_8 = _T_5 ? $signed(16'sh7f) : $signed(_T_7); // @[Mux.scala 98:16]
  wire [7:0] _T_10 = _T_8[7:0]; // @[Arithmetic.scala 126:105]
  wire [15:0] _T_13 = $signed(io_in_a) * $signed(io_in_b); // @[Arithmetic.scala 95:49]
  wire [15:0] _T_16 = $signed(_T_13) + $signed(c2); // @[Arithmetic.scala 95:54]
  wire [15:0] _T_20 = {io_in_d[7],io_in_d[7],io_in_d[7],io_in_d[7],io_in_d[7],io_in_d[7],io_in_d[7],io_in_d[7],io_in_d}; // @[Arithmetic.scala 119:61]
  wire [15:0] _T_21 = $signed(c2) >>> shift_offset; // @[PE.scala 87:23]
  wire  _T_22 = $signed(_T_21) > 16'sh7f; // @[Arithmetic.scala 126:33]
  wire  _T_23 = $signed(_T_21) < -16'sh80; // @[Arithmetic.scala 126:60]
  wire [15:0] _T_24 = _T_23 ? $signed(-16'sh80) : $signed(_T_21); // @[Mux.scala 98:16]
  wire [15:0] _T_25 = _T_22 ? $signed(16'sh7f) : $signed(_T_24); // @[Mux.scala 98:16]
  wire [7:0] _T_27 = _T_25[7:0]; // @[Arithmetic.scala 126:105]
  wire [15:0] _T_33 = $signed(_T_13) + $signed(c1); // @[Arithmetic.scala 95:54]
  wire [7:0] _GEN_1 = io_in_control_propagate ? $signed(_T_10) : $signed(_T_27); // @[PE.scala 81:30 PE.scala 82:16 PE.scala 87:16]
  wire [15:0] _GEN_22 = {{8{io_in_b[7]}},io_in_b}; // @[Arithmetic.scala 95:54]
  wire [15:0] _GEN_14 = {{8{_GEN_1[7]}},_GEN_1}; // @[PE.scala 80:95]
  assign io_out_a = io_in_a; // @[PE.scala 59:12]
  assign io_out_b = _GEN_22[7:0];
  assign io_out_c = _GEN_14[7:0];
  assign io_out_control_dataflow = io_in_control_dataflow; // @[PE.scala 60:27]
  assign io_out_control_propagate = io_in_control_propagate; // @[PE.scala 61:28]
  assign io_out_control_shift = io_in_control_shift; // @[PE.scala 62:24]
  assign io_out_id = io_in_id; // @[PE.scala 63:13]
  assign io_out_last = io_in_last; // @[PE.scala 64:15]
  assign io_out_valid = io_in_valid; // @[PE.scala 65:16]
  always @(posedge clock) begin
    if (!(~io_in_valid)) begin // @[PE.scala 109:17]
      if (io_in_control_propagate) begin // @[PE.scala 81:30]
        c1 <= _T_20; // @[PE.scala 85:10]
      end else begin
        c1 <= _T_33; // @[PE.scala 89:10]
      end
    end
    if (!(~io_in_valid)) begin // @[PE.scala 109:17]
      if (io_in_control_propagate) begin // @[PE.scala 81:30]
        c2 <= _T_16; // @[PE.scala 84:10]
      end else begin
        c2 <= _T_20; // @[PE.scala 90:10]
      end
    end
    if (io_in_valid) begin // @[Reg.scala 16:19]
      last_s <= io_in_control_propagate; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c1 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  c2 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  last_s = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tile(
  input        clock,
  input  [7:0] io_in_a_0,
  input  [7:0] io_in_a_1,
  input  [7:0] io_in_b_0,
  input  [7:0] io_in_b_1,
  input  [7:0] io_in_d_0,
  input  [7:0] io_in_d_1,
  input        io_in_control_0_dataflow,
  input        io_in_control_0_propagate,
  input  [3:0] io_in_control_0_shift,
  input        io_in_control_1_dataflow,
  input        io_in_control_1_propagate,
  input  [3:0] io_in_control_1_shift,
  input  [2:0] io_in_id_0,
  input  [2:0] io_in_id_1,
  input        io_in_last_0,
  input        io_in_last_1,
  output [7:0] io_out_a_0,
  output [7:0] io_out_a_1,
  output [7:0] io_out_c_0,
  output [7:0] io_out_c_1,
  output [7:0] io_out_b_0,
  output [7:0] io_out_b_1,
  output       io_out_control_0_dataflow,
  output       io_out_control_0_propagate,
  output [3:0] io_out_control_0_shift,
  output       io_out_control_1_dataflow,
  output       io_out_control_1_propagate,
  output [3:0] io_out_control_1_shift,
  output [2:0] io_out_id_0,
  output [2:0] io_out_id_1,
  output       io_out_last_0,
  output       io_out_last_1,
  input        io_in_valid_0,
  input        io_in_valid_1,
  output       io_out_valid_0,
  output       io_out_valid_1
);
  wire  tile_0_0_clock; // @[Tile.scala 42:44]
  wire [7:0] tile_0_0_io_in_a; // @[Tile.scala 42:44]
  wire [7:0] tile_0_0_io_in_b; // @[Tile.scala 42:44]
  wire [7:0] tile_0_0_io_in_d; // @[Tile.scala 42:44]
  wire [7:0] tile_0_0_io_out_a; // @[Tile.scala 42:44]
  wire [7:0] tile_0_0_io_out_b; // @[Tile.scala 42:44]
  wire [7:0] tile_0_0_io_out_c; // @[Tile.scala 42:44]
  wire  tile_0_0_io_in_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_0_0_io_in_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_0_0_io_in_control_shift; // @[Tile.scala 42:44]
  wire  tile_0_0_io_out_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_0_0_io_out_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_0_0_io_out_control_shift; // @[Tile.scala 42:44]
  wire [2:0] tile_0_0_io_in_id; // @[Tile.scala 42:44]
  wire [2:0] tile_0_0_io_out_id; // @[Tile.scala 42:44]
  wire  tile_0_0_io_in_last; // @[Tile.scala 42:44]
  wire  tile_0_0_io_out_last; // @[Tile.scala 42:44]
  wire  tile_0_0_io_in_valid; // @[Tile.scala 42:44]
  wire  tile_0_0_io_out_valid; // @[Tile.scala 42:44]
  wire  tile_0_1_clock; // @[Tile.scala 42:44]
  wire [7:0] tile_0_1_io_in_a; // @[Tile.scala 42:44]
  wire [7:0] tile_0_1_io_in_b; // @[Tile.scala 42:44]
  wire [7:0] tile_0_1_io_in_d; // @[Tile.scala 42:44]
  wire [7:0] tile_0_1_io_out_a; // @[Tile.scala 42:44]
  wire [7:0] tile_0_1_io_out_b; // @[Tile.scala 42:44]
  wire [7:0] tile_0_1_io_out_c; // @[Tile.scala 42:44]
  wire  tile_0_1_io_in_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_0_1_io_in_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_0_1_io_in_control_shift; // @[Tile.scala 42:44]
  wire  tile_0_1_io_out_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_0_1_io_out_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_0_1_io_out_control_shift; // @[Tile.scala 42:44]
  wire [2:0] tile_0_1_io_in_id; // @[Tile.scala 42:44]
  wire [2:0] tile_0_1_io_out_id; // @[Tile.scala 42:44]
  wire  tile_0_1_io_in_last; // @[Tile.scala 42:44]
  wire  tile_0_1_io_out_last; // @[Tile.scala 42:44]
  wire  tile_0_1_io_in_valid; // @[Tile.scala 42:44]
  wire  tile_0_1_io_out_valid; // @[Tile.scala 42:44]
  wire  tile_1_0_clock; // @[Tile.scala 42:44]
  wire [7:0] tile_1_0_io_in_a; // @[Tile.scala 42:44]
  wire [7:0] tile_1_0_io_in_b; // @[Tile.scala 42:44]
  wire [7:0] tile_1_0_io_in_d; // @[Tile.scala 42:44]
  wire [7:0] tile_1_0_io_out_a; // @[Tile.scala 42:44]
  wire [7:0] tile_1_0_io_out_b; // @[Tile.scala 42:44]
  wire [7:0] tile_1_0_io_out_c; // @[Tile.scala 42:44]
  wire  tile_1_0_io_in_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_1_0_io_in_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_1_0_io_in_control_shift; // @[Tile.scala 42:44]
  wire  tile_1_0_io_out_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_1_0_io_out_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_1_0_io_out_control_shift; // @[Tile.scala 42:44]
  wire [2:0] tile_1_0_io_in_id; // @[Tile.scala 42:44]
  wire [2:0] tile_1_0_io_out_id; // @[Tile.scala 42:44]
  wire  tile_1_0_io_in_last; // @[Tile.scala 42:44]
  wire  tile_1_0_io_out_last; // @[Tile.scala 42:44]
  wire  tile_1_0_io_in_valid; // @[Tile.scala 42:44]
  wire  tile_1_0_io_out_valid; // @[Tile.scala 42:44]
  wire  tile_1_1_clock; // @[Tile.scala 42:44]
  wire [7:0] tile_1_1_io_in_a; // @[Tile.scala 42:44]
  wire [7:0] tile_1_1_io_in_b; // @[Tile.scala 42:44]
  wire [7:0] tile_1_1_io_in_d; // @[Tile.scala 42:44]
  wire [7:0] tile_1_1_io_out_a; // @[Tile.scala 42:44]
  wire [7:0] tile_1_1_io_out_b; // @[Tile.scala 42:44]
  wire [7:0] tile_1_1_io_out_c; // @[Tile.scala 42:44]
  wire  tile_1_1_io_in_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_1_1_io_in_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_1_1_io_in_control_shift; // @[Tile.scala 42:44]
  wire  tile_1_1_io_out_control_dataflow; // @[Tile.scala 42:44]
  wire  tile_1_1_io_out_control_propagate; // @[Tile.scala 42:44]
  wire [3:0] tile_1_1_io_out_control_shift; // @[Tile.scala 42:44]
  wire [2:0] tile_1_1_io_in_id; // @[Tile.scala 42:44]
  wire [2:0] tile_1_1_io_out_id; // @[Tile.scala 42:44]
  wire  tile_1_1_io_in_last; // @[Tile.scala 42:44]
  wire  tile_1_1_io_out_last; // @[Tile.scala 42:44]
  wire  tile_1_1_io_in_valid; // @[Tile.scala 42:44]
  wire  tile_1_1_io_out_valid; // @[Tile.scala 42:44]
  PE_16 tile_0_0 ( // @[Tile.scala 42:44]
    .clock(tile_0_0_clock),
    .io_in_a(tile_0_0_io_in_a),
    .io_in_b(tile_0_0_io_in_b),
    .io_in_d(tile_0_0_io_in_d),
    .io_out_a(tile_0_0_io_out_a),
    .io_out_b(tile_0_0_io_out_b),
    .io_out_c(tile_0_0_io_out_c),
    .io_in_control_dataflow(tile_0_0_io_in_control_dataflow),
    .io_in_control_propagate(tile_0_0_io_in_control_propagate),
    .io_in_control_shift(tile_0_0_io_in_control_shift),
    .io_out_control_dataflow(tile_0_0_io_out_control_dataflow),
    .io_out_control_propagate(tile_0_0_io_out_control_propagate),
    .io_out_control_shift(tile_0_0_io_out_control_shift),
    .io_in_id(tile_0_0_io_in_id),
    .io_out_id(tile_0_0_io_out_id),
    .io_in_last(tile_0_0_io_in_last),
    .io_out_last(tile_0_0_io_out_last),
    .io_in_valid(tile_0_0_io_in_valid),
    .io_out_valid(tile_0_0_io_out_valid)
  );
  PE_16 tile_0_1 ( // @[Tile.scala 42:44]
    .clock(tile_0_1_clock),
    .io_in_a(tile_0_1_io_in_a),
    .io_in_b(tile_0_1_io_in_b),
    .io_in_d(tile_0_1_io_in_d),
    .io_out_a(tile_0_1_io_out_a),
    .io_out_b(tile_0_1_io_out_b),
    .io_out_c(tile_0_1_io_out_c),
    .io_in_control_dataflow(tile_0_1_io_in_control_dataflow),
    .io_in_control_propagate(tile_0_1_io_in_control_propagate),
    .io_in_control_shift(tile_0_1_io_in_control_shift),
    .io_out_control_dataflow(tile_0_1_io_out_control_dataflow),
    .io_out_control_propagate(tile_0_1_io_out_control_propagate),
    .io_out_control_shift(tile_0_1_io_out_control_shift),
    .io_in_id(tile_0_1_io_in_id),
    .io_out_id(tile_0_1_io_out_id),
    .io_in_last(tile_0_1_io_in_last),
    .io_out_last(tile_0_1_io_out_last),
    .io_in_valid(tile_0_1_io_in_valid),
    .io_out_valid(tile_0_1_io_out_valid)
  );
  PE_16 tile_1_0 ( // @[Tile.scala 42:44]
    .clock(tile_1_0_clock),
    .io_in_a(tile_1_0_io_in_a),
    .io_in_b(tile_1_0_io_in_b),
    .io_in_d(tile_1_0_io_in_d),
    .io_out_a(tile_1_0_io_out_a),
    .io_out_b(tile_1_0_io_out_b),
    .io_out_c(tile_1_0_io_out_c),
    .io_in_control_dataflow(tile_1_0_io_in_control_dataflow),
    .io_in_control_propagate(tile_1_0_io_in_control_propagate),
    .io_in_control_shift(tile_1_0_io_in_control_shift),
    .io_out_control_dataflow(tile_1_0_io_out_control_dataflow),
    .io_out_control_propagate(tile_1_0_io_out_control_propagate),
    .io_out_control_shift(tile_1_0_io_out_control_shift),
    .io_in_id(tile_1_0_io_in_id),
    .io_out_id(tile_1_0_io_out_id),
    .io_in_last(tile_1_0_io_in_last),
    .io_out_last(tile_1_0_io_out_last),
    .io_in_valid(tile_1_0_io_in_valid),
    .io_out_valid(tile_1_0_io_out_valid)
  );
  PE_16 tile_1_1 ( // @[Tile.scala 42:44]
    .clock(tile_1_1_clock),
    .io_in_a(tile_1_1_io_in_a),
    .io_in_b(tile_1_1_io_in_b),
    .io_in_d(tile_1_1_io_in_d),
    .io_out_a(tile_1_1_io_out_a),
    .io_out_b(tile_1_1_io_out_b),
    .io_out_c(tile_1_1_io_out_c),
    .io_in_control_dataflow(tile_1_1_io_in_control_dataflow),
    .io_in_control_propagate(tile_1_1_io_in_control_propagate),
    .io_in_control_shift(tile_1_1_io_in_control_shift),
    .io_out_control_dataflow(tile_1_1_io_out_control_dataflow),
    .io_out_control_propagate(tile_1_1_io_out_control_propagate),
    .io_out_control_shift(tile_1_1_io_out_control_shift),
    .io_in_id(tile_1_1_io_in_id),
    .io_out_id(tile_1_1_io_out_id),
    .io_in_last(tile_1_1_io_in_last),
    .io_out_last(tile_1_1_io_out_last),
    .io_in_valid(tile_1_1_io_in_valid),
    .io_out_valid(tile_1_1_io_out_valid)
  );
  assign io_out_a_0 = tile_0_1_io_out_a; // @[Tile.scala 123:17]
  assign io_out_a_1 = tile_1_1_io_out_a; // @[Tile.scala 123:17]
  assign io_out_c_0 = tile_1_0_io_out_c; // @[Tile.scala 111:17]
  assign io_out_c_1 = tile_1_1_io_out_c; // @[Tile.scala 111:17]
  assign io_out_b_0 = tile_1_0_io_out_b; // @[Tile.scala 116:17]
  assign io_out_b_1 = tile_1_1_io_out_b; // @[Tile.scala 116:17]
  assign io_out_control_0_dataflow = tile_1_0_io_out_control_dataflow; // @[Tile.scala 112:23]
  assign io_out_control_0_propagate = tile_1_0_io_out_control_propagate; // @[Tile.scala 112:23]
  assign io_out_control_0_shift = tile_1_0_io_out_control_shift; // @[Tile.scala 112:23]
  assign io_out_control_1_dataflow = tile_1_1_io_out_control_dataflow; // @[Tile.scala 112:23]
  assign io_out_control_1_propagate = tile_1_1_io_out_control_propagate; // @[Tile.scala 112:23]
  assign io_out_control_1_shift = tile_1_1_io_out_control_shift; // @[Tile.scala 112:23]
  assign io_out_id_0 = tile_1_0_io_out_id; // @[Tile.scala 113:18]
  assign io_out_id_1 = tile_1_1_io_out_id; // @[Tile.scala 113:18]
  assign io_out_last_0 = tile_1_0_io_out_last; // @[Tile.scala 114:20]
  assign io_out_last_1 = tile_1_1_io_out_last; // @[Tile.scala 114:20]
  assign io_out_valid_0 = tile_1_0_io_out_valid; // @[Tile.scala 115:21]
  assign io_out_valid_1 = tile_1_1_io_out_valid; // @[Tile.scala 115:21]
  assign tile_0_0_clock = clock;
  assign tile_0_0_io_in_a = io_in_a_0; // @[Tile.scala 50:20]
  assign tile_0_0_io_in_b = io_in_b_0; // @[Tile.scala 59:20]
  assign tile_0_0_io_in_d = io_in_d_0; // @[Tile.scala 68:20]
  assign tile_0_0_io_in_control_dataflow = io_in_control_0_dataflow; // @[Tile.scala 77:26]
  assign tile_0_0_io_in_control_propagate = io_in_control_0_propagate; // @[Tile.scala 77:26]
  assign tile_0_0_io_in_control_shift = io_in_control_0_shift; // @[Tile.scala 77:26]
  assign tile_0_0_io_in_id = io_in_id_0; // @[Tile.scala 95:21]
  assign tile_0_0_io_in_last = io_in_last_0; // @[Tile.scala 104:23]
  assign tile_0_0_io_in_valid = io_in_valid_0; // @[Tile.scala 86:24]
  assign tile_0_1_clock = clock;
  assign tile_0_1_io_in_a = tile_0_0_io_out_a; // @[Tile.scala 50:20]
  assign tile_0_1_io_in_b = io_in_b_1; // @[Tile.scala 59:20]
  assign tile_0_1_io_in_d = io_in_d_1; // @[Tile.scala 68:20]
  assign tile_0_1_io_in_control_dataflow = io_in_control_1_dataflow; // @[Tile.scala 77:26]
  assign tile_0_1_io_in_control_propagate = io_in_control_1_propagate; // @[Tile.scala 77:26]
  assign tile_0_1_io_in_control_shift = io_in_control_1_shift; // @[Tile.scala 77:26]
  assign tile_0_1_io_in_id = io_in_id_1; // @[Tile.scala 95:21]
  assign tile_0_1_io_in_last = io_in_last_1; // @[Tile.scala 104:23]
  assign tile_0_1_io_in_valid = io_in_valid_1; // @[Tile.scala 86:24]
  assign tile_1_0_clock = clock;
  assign tile_1_0_io_in_a = io_in_a_1; // @[Tile.scala 50:20]
  assign tile_1_0_io_in_b = tile_0_0_io_out_b; // @[Tile.scala 59:20]
  assign tile_1_0_io_in_d = tile_0_0_io_out_c; // @[Tile.scala 68:20]
  assign tile_1_0_io_in_control_dataflow = tile_0_0_io_out_control_dataflow; // @[Tile.scala 77:26]
  assign tile_1_0_io_in_control_propagate = tile_0_0_io_out_control_propagate; // @[Tile.scala 77:26]
  assign tile_1_0_io_in_control_shift = tile_0_0_io_out_control_shift; // @[Tile.scala 77:26]
  assign tile_1_0_io_in_id = tile_0_0_io_out_id; // @[Tile.scala 95:21]
  assign tile_1_0_io_in_last = tile_0_0_io_out_last; // @[Tile.scala 104:23]
  assign tile_1_0_io_in_valid = tile_0_0_io_out_valid; // @[Tile.scala 86:24]
  assign tile_1_1_clock = clock;
  assign tile_1_1_io_in_a = tile_1_0_io_out_a; // @[Tile.scala 50:20]
  assign tile_1_1_io_in_b = tile_0_1_io_out_b; // @[Tile.scala 59:20]
  assign tile_1_1_io_in_d = tile_0_1_io_out_c; // @[Tile.scala 68:20]
  assign tile_1_1_io_in_control_dataflow = tile_0_1_io_out_control_dataflow; // @[Tile.scala 77:26]
  assign tile_1_1_io_in_control_propagate = tile_0_1_io_out_control_propagate; // @[Tile.scala 77:26]
  assign tile_1_1_io_in_control_shift = tile_0_1_io_out_control_shift; // @[Tile.scala 77:26]
  assign tile_1_1_io_in_id = tile_0_1_io_out_id; // @[Tile.scala 95:21]
  assign tile_1_1_io_in_last = tile_0_1_io_out_last; // @[Tile.scala 104:23]
  assign tile_1_1_io_in_valid = tile_0_1_io_out_valid; // @[Tile.scala 86:24]
endmodule
module Mesh(
  input        clock,
  input  [7:0] io_in_a_0_0,
  input  [7:0] io_in_a_0_1,
  input  [7:0] io_in_a_1_0,
  input  [7:0] io_in_a_1_1,
  input  [7:0] io_in_b_0_0,
  input  [7:0] io_in_b_0_1,
  input  [7:0] io_in_b_1_0,
  input  [7:0] io_in_b_1_1,
  input  [7:0] io_in_d_0_0,
  input  [7:0] io_in_d_0_1,
  input  [7:0] io_in_d_1_0,
  input  [7:0] io_in_d_1_1,
  input        io_in_control_0_0_dataflow,
  input        io_in_control_0_0_propagate,
  input  [3:0] io_in_control_0_0_shift,
  input        io_in_control_0_1_dataflow,
  input        io_in_control_0_1_propagate,
  input  [3:0] io_in_control_0_1_shift,
  input        io_in_control_1_0_dataflow,
  input        io_in_control_1_0_propagate,
  input  [3:0] io_in_control_1_0_shift,
  input        io_in_control_1_1_dataflow,
  input        io_in_control_1_1_propagate,
  input  [3:0] io_in_control_1_1_shift,
  input  [2:0] io_in_id_0_0,
  input  [2:0] io_in_id_0_1,
  input  [2:0] io_in_id_1_0,
  input  [2:0] io_in_id_1_1,
  input        io_in_last_0_0,
  input        io_in_last_0_1,
  input        io_in_last_1_0,
  input        io_in_last_1_1,
  output [7:0] io_out_b_0_0,
  output [7:0] io_out_b_0_1,
  output [7:0] io_out_b_1_0,
  output [7:0] io_out_b_1_1,
  output [7:0] io_out_c_0_0,
  output [7:0] io_out_c_0_1,
  output [7:0] io_out_c_1_0,
  output [7:0] io_out_c_1_1,
  input        io_in_valid_0_0,
  input        io_in_valid_0_1,
  input        io_in_valid_1_0,
  input        io_in_valid_1_1,
  output       io_out_valid_0_0,
  output       io_out_control_0_0_dataflow,
  output [2:0] io_out_id_0_0,
  output       io_out_last_0_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
`endif // RANDOMIZE_REG_INIT
  wire  mesh_0_0_clock; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_in_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_in_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_in_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_in_b_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_in_d_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_in_d_1; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_0_io_in_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_0_io_in_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_0_io_in_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_0_io_in_id_1; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_last_0; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_last_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_out_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_out_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_out_c_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_out_c_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_out_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_0_io_out_b_1; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_0_io_out_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_0_io_out_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_0_io_out_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_0_io_out_id_1; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_last_0; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_last_1; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_in_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_0_0_io_out_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_clock; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_in_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_in_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_in_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_in_b_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_in_d_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_in_d_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_1_io_in_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_1_io_in_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_1_io_in_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_1_io_in_id_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_last_0; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_last_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_out_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_out_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_out_c_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_out_c_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_out_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_0_1_io_out_b_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_1_io_out_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_0_1_io_out_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_1_io_out_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_0_1_io_out_id_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_last_0; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_last_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_in_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_0_1_io_out_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_clock; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_in_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_in_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_in_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_in_b_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_in_d_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_in_d_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_0_io_in_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_0_io_in_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_0_io_in_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_0_io_in_id_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_last_0; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_last_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_out_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_out_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_out_c_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_out_c_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_out_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_0_io_out_b_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_0_io_out_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_0_io_out_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_0_io_out_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_0_io_out_id_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_last_0; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_last_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_in_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_1_0_io_out_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_clock; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_in_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_in_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_in_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_in_b_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_in_d_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_in_d_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_1_io_in_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_1_io_in_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_1_io_in_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_1_io_in_id_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_last_0; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_last_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_out_a_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_out_a_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_out_c_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_out_c_1; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_out_b_0; // @[Mesh.scala 38:68]
  wire [7:0] mesh_1_1_io_out_b_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_control_0_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_control_0_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_1_io_out_control_0_shift; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_control_1_dataflow; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_control_1_propagate; // @[Mesh.scala 38:68]
  wire [3:0] mesh_1_1_io_out_control_1_shift; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_1_io_out_id_0; // @[Mesh.scala 38:68]
  wire [2:0] mesh_1_1_io_out_id_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_last_0; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_last_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_in_valid_1; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_valid_0; // @[Mesh.scala 38:68]
  wire  mesh_1_1_io_out_valid_1; // @[Mesh.scala 38:68]
  reg [7:0] r__0; // @[Reg.scala 15:16]
  reg [7:0] r__1; // @[Reg.scala 15:16]
  reg [7:0] r_1_0; // @[Reg.scala 15:16]
  reg [7:0] r_1_1; // @[Reg.scala 15:16]
  reg [7:0] r_2_0; // @[Reg.scala 15:16]
  reg [7:0] r_2_1; // @[Reg.scala 15:16]
  reg [7:0] r_3_0; // @[Reg.scala 15:16]
  reg [7:0] r_3_1; // @[Reg.scala 15:16]
  reg [7:0] r_4_0; // @[Reg.scala 15:16]
  reg [7:0] r_4_1; // @[Reg.scala 15:16]
  reg [7:0] r_5_0; // @[Reg.scala 15:16]
  reg [7:0] r_5_1; // @[Reg.scala 15:16]
  reg [7:0] r_6_0; // @[Reg.scala 15:16]
  reg [7:0] r_6_1; // @[Reg.scala 15:16]
  reg [7:0] r_7_0; // @[Reg.scala 15:16]
  reg [7:0] r_7_1; // @[Reg.scala 15:16]
  reg  v; // @[Valid.scala 117:22]
  reg [7:0] b__0; // @[Reg.scala 15:16]
  reg [7:0] b__1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits__0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits__1; // @[Reg.scala 15:16]
  reg  v_1; // @[Valid.scala 117:22]
  reg [7:0] b_1_0; // @[Reg.scala 15:16]
  reg [7:0] b_1_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_1_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_1_1; // @[Reg.scala 15:16]
  reg  v_2; // @[Valid.scala 117:22]
  reg [7:0] b_2_0; // @[Reg.scala 15:16]
  reg [7:0] b_2_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_2_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_2_1; // @[Reg.scala 15:16]
  reg  v_3; // @[Valid.scala 117:22]
  reg [7:0] b_3_0; // @[Reg.scala 15:16]
  reg [7:0] b_3_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_3_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_3_1; // @[Reg.scala 15:16]
  reg  v_4; // @[Valid.scala 117:22]
  reg [7:0] b_4_0; // @[Reg.scala 15:16]
  reg [7:0] b_4_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_4_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_4_1; // @[Reg.scala 15:16]
  reg  v_5; // @[Valid.scala 117:22]
  reg [7:0] b_5_0; // @[Reg.scala 15:16]
  reg [7:0] b_5_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_5_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_5_1; // @[Reg.scala 15:16]
  reg  v_6; // @[Valid.scala 117:22]
  reg [7:0] b_6_0; // @[Reg.scala 15:16]
  reg [7:0] b_6_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_6_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_6_1; // @[Reg.scala 15:16]
  reg  v_7; // @[Valid.scala 117:22]
  reg [7:0] b_7_0; // @[Reg.scala 15:16]
  reg [7:0] b_7_1; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_7_0; // @[Reg.scala 15:16]
  reg [7:0] outPipe_bits_7_1; // @[Reg.scala 15:16]
  reg  v_8; // @[Valid.scala 117:22]
  reg [3:0] b_8; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_8; // @[Reg.scala 15:16]
  reg  v_9; // @[Valid.scala 117:22]
  reg  b_9; // @[Reg.scala 15:16]
  reg  outPipe_bits_9; // @[Reg.scala 15:16]
  reg  v_10; // @[Valid.scala 117:22]
  reg  b_10; // @[Reg.scala 15:16]
  reg  outPipe_bits_10; // @[Reg.scala 15:16]
  reg  v_11; // @[Valid.scala 117:22]
  reg [3:0] b_11; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_11; // @[Reg.scala 15:16]
  reg  v_12; // @[Valid.scala 117:22]
  reg  b_12; // @[Reg.scala 15:16]
  reg  outPipe_bits_12; // @[Reg.scala 15:16]
  reg  v_13; // @[Valid.scala 117:22]
  reg  b_13; // @[Reg.scala 15:16]
  reg  outPipe_bits_13; // @[Reg.scala 15:16]
  reg  v_14; // @[Valid.scala 117:22]
  reg [3:0] b_14; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_14; // @[Reg.scala 15:16]
  reg  v_15; // @[Valid.scala 117:22]
  reg  b_15; // @[Reg.scala 15:16]
  reg  outPipe_bits_15; // @[Reg.scala 15:16]
  reg  v_16; // @[Valid.scala 117:22]
  reg  b_16; // @[Reg.scala 15:16]
  reg  outPipe_bits_16; // @[Reg.scala 15:16]
  reg  v_17; // @[Valid.scala 117:22]
  reg [3:0] b_17; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_17; // @[Reg.scala 15:16]
  reg  v_18; // @[Valid.scala 117:22]
  reg  b_18; // @[Reg.scala 15:16]
  reg  outPipe_bits_18; // @[Reg.scala 15:16]
  reg  v_19; // @[Valid.scala 117:22]
  reg  b_19; // @[Reg.scala 15:16]
  reg  outPipe_bits_19; // @[Reg.scala 15:16]
  reg  v_20; // @[Valid.scala 117:22]
  reg [3:0] b_20; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_20; // @[Reg.scala 15:16]
  reg  v_21; // @[Valid.scala 117:22]
  reg  b_21; // @[Reg.scala 15:16]
  reg  outPipe_bits_21; // @[Reg.scala 15:16]
  reg  v_22; // @[Valid.scala 117:22]
  reg  b_22; // @[Reg.scala 15:16]
  reg  outPipe_bits_22; // @[Reg.scala 15:16]
  reg  v_23; // @[Valid.scala 117:22]
  reg [3:0] b_23; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_23; // @[Reg.scala 15:16]
  reg  v_24; // @[Valid.scala 117:22]
  reg  b_24; // @[Reg.scala 15:16]
  reg  outPipe_bits_24; // @[Reg.scala 15:16]
  reg  v_25; // @[Valid.scala 117:22]
  reg  b_25; // @[Reg.scala 15:16]
  reg  outPipe_bits_25; // @[Reg.scala 15:16]
  reg  v_26; // @[Valid.scala 117:22]
  reg [3:0] b_26; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_26; // @[Reg.scala 15:16]
  reg  v_27; // @[Valid.scala 117:22]
  reg  b_27; // @[Reg.scala 15:16]
  reg  outPipe_bits_27; // @[Reg.scala 15:16]
  reg  v_28; // @[Valid.scala 117:22]
  reg  b_28; // @[Reg.scala 15:16]
  reg  outPipe_bits_28; // @[Reg.scala 15:16]
  reg  v_29; // @[Valid.scala 117:22]
  reg [3:0] b_29; // @[Reg.scala 15:16]
  reg [3:0] outPipe_bits_29; // @[Reg.scala 15:16]
  reg  v_30; // @[Valid.scala 117:22]
  reg  b_30; // @[Reg.scala 15:16]
  reg  outPipe_bits_30; // @[Reg.scala 15:16]
  reg  v_31; // @[Valid.scala 117:22]
  reg  b_31; // @[Reg.scala 15:16]
  reg  outPipe_bits_31; // @[Reg.scala 15:16]
  reg  r_8_0; // @[Reg.scala 15:16]
  reg  r_8_1; // @[Reg.scala 15:16]
  reg  r_9_0; // @[Reg.scala 15:16]
  reg  r_9_1; // @[Reg.scala 15:16]
  reg  r_10_0; // @[Reg.scala 15:16]
  reg  r_10_1; // @[Reg.scala 15:16]
  reg  r_11_0; // @[Reg.scala 15:16]
  reg  r_11_1; // @[Reg.scala 15:16]
  reg  r_12_0; // @[Reg.scala 15:16]
  reg  r_12_1; // @[Reg.scala 15:16]
  reg  r_13_0; // @[Reg.scala 15:16]
  reg  r_13_1; // @[Reg.scala 15:16]
  reg  r_14_0; // @[Reg.scala 15:16]
  reg  r_14_1; // @[Reg.scala 15:16]
  reg  r_15_0; // @[Reg.scala 15:16]
  reg  r_15_1; // @[Reg.scala 15:16]
  reg [2:0] r_16_0; // @[Reg.scala 15:16]
  reg [2:0] r_16_1; // @[Reg.scala 15:16]
  reg [2:0] r_17_0; // @[Reg.scala 15:16]
  reg [2:0] r_17_1; // @[Reg.scala 15:16]
  reg [2:0] r_18_0; // @[Reg.scala 15:16]
  reg [2:0] r_18_1; // @[Reg.scala 15:16]
  reg [2:0] r_19_0; // @[Reg.scala 15:16]
  reg [2:0] r_19_1; // @[Reg.scala 15:16]
  reg [2:0] r_20_0; // @[Reg.scala 15:16]
  reg [2:0] r_20_1; // @[Reg.scala 15:16]
  reg [2:0] r_21_0; // @[Reg.scala 15:16]
  reg [2:0] r_21_1; // @[Reg.scala 15:16]
  reg [2:0] r_22_0; // @[Reg.scala 15:16]
  reg [2:0] r_22_1; // @[Reg.scala 15:16]
  reg [2:0] r_23_0; // @[Reg.scala 15:16]
  reg [2:0] r_23_1; // @[Reg.scala 15:16]
  reg  r_24_0; // @[Reg.scala 15:16]
  reg  r_24_1; // @[Reg.scala 15:16]
  reg  r_25_0; // @[Reg.scala 15:16]
  reg  r_25_1; // @[Reg.scala 15:16]
  reg  r_26_0; // @[Reg.scala 15:16]
  reg  r_26_1; // @[Reg.scala 15:16]
  reg  r_27_0; // @[Reg.scala 15:16]
  reg  r_27_1; // @[Reg.scala 15:16]
  reg  r_28_0; // @[Reg.scala 15:16]
  reg  r_28_1; // @[Reg.scala 15:16]
  reg  r_29_0; // @[Reg.scala 15:16]
  reg  r_29_1; // @[Reg.scala 15:16]
  reg  r_30_0; // @[Reg.scala 15:16]
  reg  r_30_1; // @[Reg.scala 15:16]
  reg  r_31_0; // @[Reg.scala 15:16]
  reg  r_31_1; // @[Reg.scala 15:16]
  reg [7:0] r_32_0; // @[Reg.scala 15:16]
  reg [7:0] r_32_1; // @[Reg.scala 15:16]
  reg [7:0] r_33_0; // @[Reg.scala 15:16]
  reg [7:0] r_33_1; // @[Reg.scala 15:16]
  reg  r_34_0; // @[Reg.scala 15:16]
  reg  r_35_0_dataflow; // @[Reg.scala 15:16]
  reg [2:0] r_36_0; // @[Reg.scala 15:16]
  reg  r_37_0; // @[Reg.scala 15:16]
  reg [7:0] r_38_0; // @[Reg.scala 15:16]
  reg [7:0] r_38_1; // @[Reg.scala 15:16]
  reg [7:0] r_39_0; // @[Reg.scala 15:16]
  reg [7:0] r_39_1; // @[Reg.scala 15:16]
  Tile mesh_0_0 ( // @[Mesh.scala 38:68]
    .clock(mesh_0_0_clock),
    .io_in_a_0(mesh_0_0_io_in_a_0),
    .io_in_a_1(mesh_0_0_io_in_a_1),
    .io_in_b_0(mesh_0_0_io_in_b_0),
    .io_in_b_1(mesh_0_0_io_in_b_1),
    .io_in_d_0(mesh_0_0_io_in_d_0),
    .io_in_d_1(mesh_0_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_0_io_in_control_1_shift),
    .io_in_id_0(mesh_0_0_io_in_id_0),
    .io_in_id_1(mesh_0_0_io_in_id_1),
    .io_in_last_0(mesh_0_0_io_in_last_0),
    .io_in_last_1(mesh_0_0_io_in_last_1),
    .io_out_a_0(mesh_0_0_io_out_a_0),
    .io_out_a_1(mesh_0_0_io_out_a_1),
    .io_out_c_0(mesh_0_0_io_out_c_0),
    .io_out_c_1(mesh_0_0_io_out_c_1),
    .io_out_b_0(mesh_0_0_io_out_b_0),
    .io_out_b_1(mesh_0_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_0_io_out_control_1_shift),
    .io_out_id_0(mesh_0_0_io_out_id_0),
    .io_out_id_1(mesh_0_0_io_out_id_1),
    .io_out_last_0(mesh_0_0_io_out_last_0),
    .io_out_last_1(mesh_0_0_io_out_last_1),
    .io_in_valid_0(mesh_0_0_io_in_valid_0),
    .io_in_valid_1(mesh_0_0_io_in_valid_1),
    .io_out_valid_0(mesh_0_0_io_out_valid_0),
    .io_out_valid_1(mesh_0_0_io_out_valid_1)
  );
  Tile mesh_0_1 ( // @[Mesh.scala 38:68]
    .clock(mesh_0_1_clock),
    .io_in_a_0(mesh_0_1_io_in_a_0),
    .io_in_a_1(mesh_0_1_io_in_a_1),
    .io_in_b_0(mesh_0_1_io_in_b_0),
    .io_in_b_1(mesh_0_1_io_in_b_1),
    .io_in_d_0(mesh_0_1_io_in_d_0),
    .io_in_d_1(mesh_0_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_0_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_0_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_0_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_0_1_io_in_control_1_shift),
    .io_in_id_0(mesh_0_1_io_in_id_0),
    .io_in_id_1(mesh_0_1_io_in_id_1),
    .io_in_last_0(mesh_0_1_io_in_last_0),
    .io_in_last_1(mesh_0_1_io_in_last_1),
    .io_out_a_0(mesh_0_1_io_out_a_0),
    .io_out_a_1(mesh_0_1_io_out_a_1),
    .io_out_c_0(mesh_0_1_io_out_c_0),
    .io_out_c_1(mesh_0_1_io_out_c_1),
    .io_out_b_0(mesh_0_1_io_out_b_0),
    .io_out_b_1(mesh_0_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_0_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_0_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_0_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_0_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_0_1_io_out_control_1_shift),
    .io_out_id_0(mesh_0_1_io_out_id_0),
    .io_out_id_1(mesh_0_1_io_out_id_1),
    .io_out_last_0(mesh_0_1_io_out_last_0),
    .io_out_last_1(mesh_0_1_io_out_last_1),
    .io_in_valid_0(mesh_0_1_io_in_valid_0),
    .io_in_valid_1(mesh_0_1_io_in_valid_1),
    .io_out_valid_0(mesh_0_1_io_out_valid_0),
    .io_out_valid_1(mesh_0_1_io_out_valid_1)
  );
  Tile mesh_1_0 ( // @[Mesh.scala 38:68]
    .clock(mesh_1_0_clock),
    .io_in_a_0(mesh_1_0_io_in_a_0),
    .io_in_a_1(mesh_1_0_io_in_a_1),
    .io_in_b_0(mesh_1_0_io_in_b_0),
    .io_in_b_1(mesh_1_0_io_in_b_1),
    .io_in_d_0(mesh_1_0_io_in_d_0),
    .io_in_d_1(mesh_1_0_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_0_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_0_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_0_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_0_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_0_io_in_control_1_shift),
    .io_in_id_0(mesh_1_0_io_in_id_0),
    .io_in_id_1(mesh_1_0_io_in_id_1),
    .io_in_last_0(mesh_1_0_io_in_last_0),
    .io_in_last_1(mesh_1_0_io_in_last_1),
    .io_out_a_0(mesh_1_0_io_out_a_0),
    .io_out_a_1(mesh_1_0_io_out_a_1),
    .io_out_c_0(mesh_1_0_io_out_c_0),
    .io_out_c_1(mesh_1_0_io_out_c_1),
    .io_out_b_0(mesh_1_0_io_out_b_0),
    .io_out_b_1(mesh_1_0_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_0_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_0_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_0_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_0_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_0_io_out_control_1_shift),
    .io_out_id_0(mesh_1_0_io_out_id_0),
    .io_out_id_1(mesh_1_0_io_out_id_1),
    .io_out_last_0(mesh_1_0_io_out_last_0),
    .io_out_last_1(mesh_1_0_io_out_last_1),
    .io_in_valid_0(mesh_1_0_io_in_valid_0),
    .io_in_valid_1(mesh_1_0_io_in_valid_1),
    .io_out_valid_0(mesh_1_0_io_out_valid_0),
    .io_out_valid_1(mesh_1_0_io_out_valid_1)
  );
  Tile mesh_1_1 ( // @[Mesh.scala 38:68]
    .clock(mesh_1_1_clock),
    .io_in_a_0(mesh_1_1_io_in_a_0),
    .io_in_a_1(mesh_1_1_io_in_a_1),
    .io_in_b_0(mesh_1_1_io_in_b_0),
    .io_in_b_1(mesh_1_1_io_in_b_1),
    .io_in_d_0(mesh_1_1_io_in_d_0),
    .io_in_d_1(mesh_1_1_io_in_d_1),
    .io_in_control_0_dataflow(mesh_1_1_io_in_control_0_dataflow),
    .io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_1_io_in_control_0_shift),
    .io_in_control_1_dataflow(mesh_1_1_io_in_control_1_dataflow),
    .io_in_control_1_propagate(mesh_1_1_io_in_control_1_propagate),
    .io_in_control_1_shift(mesh_1_1_io_in_control_1_shift),
    .io_in_id_0(mesh_1_1_io_in_id_0),
    .io_in_id_1(mesh_1_1_io_in_id_1),
    .io_in_last_0(mesh_1_1_io_in_last_0),
    .io_in_last_1(mesh_1_1_io_in_last_1),
    .io_out_a_0(mesh_1_1_io_out_a_0),
    .io_out_a_1(mesh_1_1_io_out_a_1),
    .io_out_c_0(mesh_1_1_io_out_c_0),
    .io_out_c_1(mesh_1_1_io_out_c_1),
    .io_out_b_0(mesh_1_1_io_out_b_0),
    .io_out_b_1(mesh_1_1_io_out_b_1),
    .io_out_control_0_dataflow(mesh_1_1_io_out_control_0_dataflow),
    .io_out_control_0_propagate(mesh_1_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_1_io_out_control_0_shift),
    .io_out_control_1_dataflow(mesh_1_1_io_out_control_1_dataflow),
    .io_out_control_1_propagate(mesh_1_1_io_out_control_1_propagate),
    .io_out_control_1_shift(mesh_1_1_io_out_control_1_shift),
    .io_out_id_0(mesh_1_1_io_out_id_0),
    .io_out_id_1(mesh_1_1_io_out_id_1),
    .io_out_last_0(mesh_1_1_io_out_last_0),
    .io_out_last_1(mesh_1_1_io_out_last_1),
    .io_in_valid_0(mesh_1_1_io_in_valid_0),
    .io_in_valid_1(mesh_1_1_io_in_valid_1),
    .io_out_valid_0(mesh_1_1_io_out_valid_0),
    .io_out_valid_1(mesh_1_1_io_out_valid_1)
  );
  assign io_out_b_0_0 = r_32_0; // @[Mesh.scala 121:7]
  assign io_out_b_0_1 = r_32_1; // @[Mesh.scala 121:7]
  assign io_out_b_1_0 = r_38_0; // @[Mesh.scala 121:7]
  assign io_out_b_1_1 = r_38_1; // @[Mesh.scala 121:7]
  assign io_out_c_0_0 = r_33_0; // @[Mesh.scala 122:7]
  assign io_out_c_0_1 = r_33_1; // @[Mesh.scala 122:7]
  assign io_out_c_1_0 = r_39_0; // @[Mesh.scala 122:7]
  assign io_out_c_1_1 = r_39_1; // @[Mesh.scala 122:7]
  assign io_out_valid_0_0 = r_34_0; // @[Mesh.scala 123:7]
  assign io_out_control_0_0_dataflow = r_35_0_dataflow; // @[Mesh.scala 124:10]
  assign io_out_id_0_0 = r_36_0; // @[Mesh.scala 125:8]
  assign io_out_last_0_0 = r_37_0; // @[Mesh.scala 126:10]
  assign mesh_0_0_clock = clock;
  assign mesh_0_0_io_in_a_0 = r_1_0; // @[Mesh.scala 52:22]
  assign mesh_0_0_io_in_a_1 = r_1_1; // @[Mesh.scala 52:22]
  assign mesh_0_0_io_in_b_0 = outPipe_bits__0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_b_1 = outPipe_bits__1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_d_0 = outPipe_bits_4_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_d_1 = outPipe_bits_4_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_control_0_dataflow = outPipe_bits_9; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_control_0_propagate = outPipe_bits_10; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_control_0_shift = outPipe_bits_8; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_control_1_dataflow = outPipe_bits_12; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_control_1_propagate = outPipe_bits_13; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_control_1_shift = outPipe_bits_11; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_0_io_in_id_0 = r_17_0; // @[Mesh.scala 102:23]
  assign mesh_0_0_io_in_id_1 = r_17_1; // @[Mesh.scala 102:23]
  assign mesh_0_0_io_in_last_0 = r_25_0; // @[Mesh.scala 111:25]
  assign mesh_0_0_io_in_last_1 = r_25_1; // @[Mesh.scala 111:25]
  assign mesh_0_0_io_in_valid_0 = r_9_0; // @[Mesh.scala 93:26]
  assign mesh_0_0_io_in_valid_1 = r_9_1; // @[Mesh.scala 93:26]
  assign mesh_0_1_clock = clock;
  assign mesh_0_1_io_in_a_0 = r_3_0; // @[Mesh.scala 52:22]
  assign mesh_0_1_io_in_a_1 = r_3_1; // @[Mesh.scala 52:22]
  assign mesh_0_1_io_in_b_0 = outPipe_bits_2_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_b_1 = outPipe_bits_2_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_d_0 = outPipe_bits_6_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_d_1 = outPipe_bits_6_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_control_0_dataflow = outPipe_bits_21; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_control_0_propagate = outPipe_bits_22; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_control_0_shift = outPipe_bits_20; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_control_1_dataflow = outPipe_bits_24; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_control_1_propagate = outPipe_bits_25; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_control_1_shift = outPipe_bits_23; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_0_1_io_in_id_0 = r_21_0; // @[Mesh.scala 102:23]
  assign mesh_0_1_io_in_id_1 = r_21_1; // @[Mesh.scala 102:23]
  assign mesh_0_1_io_in_last_0 = r_29_0; // @[Mesh.scala 111:25]
  assign mesh_0_1_io_in_last_1 = r_29_1; // @[Mesh.scala 111:25]
  assign mesh_0_1_io_in_valid_0 = r_13_0; // @[Mesh.scala 93:26]
  assign mesh_0_1_io_in_valid_1 = r_13_1; // @[Mesh.scala 93:26]
  assign mesh_1_0_clock = clock;
  assign mesh_1_0_io_in_a_0 = r_5_0; // @[Mesh.scala 52:22]
  assign mesh_1_0_io_in_a_1 = r_5_1; // @[Mesh.scala 52:22]
  assign mesh_1_0_io_in_b_0 = outPipe_bits_1_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_b_1 = outPipe_bits_1_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_d_0 = outPipe_bits_5_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_d_1 = outPipe_bits_5_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_control_0_dataflow = outPipe_bits_15; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_control_0_propagate = outPipe_bits_16; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_control_0_shift = outPipe_bits_14; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_control_1_dataflow = outPipe_bits_18; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_control_1_propagate = outPipe_bits_19; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_control_1_shift = outPipe_bits_17; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_0_io_in_id_0 = r_19_0; // @[Mesh.scala 102:23]
  assign mesh_1_0_io_in_id_1 = r_19_1; // @[Mesh.scala 102:23]
  assign mesh_1_0_io_in_last_0 = r_27_0; // @[Mesh.scala 111:25]
  assign mesh_1_0_io_in_last_1 = r_27_1; // @[Mesh.scala 111:25]
  assign mesh_1_0_io_in_valid_0 = r_11_0; // @[Mesh.scala 93:26]
  assign mesh_1_0_io_in_valid_1 = r_11_1; // @[Mesh.scala 93:26]
  assign mesh_1_1_clock = clock;
  assign mesh_1_1_io_in_a_0 = r_7_0; // @[Mesh.scala 52:22]
  assign mesh_1_1_io_in_a_1 = r_7_1; // @[Mesh.scala 52:22]
  assign mesh_1_1_io_in_b_0 = outPipe_bits_3_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_b_1 = outPipe_bits_3_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_d_0 = outPipe_bits_7_0; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_d_1 = outPipe_bits_7_1; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_control_0_dataflow = outPipe_bits_27; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_control_0_propagate = outPipe_bits_28; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_control_0_shift = outPipe_bits_26; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_control_1_dataflow = outPipe_bits_30; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_control_1_propagate = outPipe_bits_31; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_control_1_shift = outPipe_bits_29; // @[Valid.scala 112:21 Valid.scala 114:16]
  assign mesh_1_1_io_in_id_0 = r_23_0; // @[Mesh.scala 102:23]
  assign mesh_1_1_io_in_id_1 = r_23_1; // @[Mesh.scala 102:23]
  assign mesh_1_1_io_in_last_0 = r_31_0; // @[Mesh.scala 111:25]
  assign mesh_1_1_io_in_last_1 = r_31_1; // @[Mesh.scala 111:25]
  assign mesh_1_1_io_in_valid_0 = r_15_0; // @[Mesh.scala 93:26]
  assign mesh_1_1_io_in_valid_1 = r_15_1; // @[Mesh.scala 93:26]
  always @(posedge clock) begin
    r__0 <= io_in_a_0_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r__1 <= io_in_a_0_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_1_0 <= r__0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_1_1 <= r__1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_2_0 <= mesh_0_0_io_out_a_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_2_1 <= mesh_0_0_io_out_a_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_3_0 <= r_2_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_3_1 <= r_2_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_4_0 <= io_in_a_1_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_4_1 <= io_in_a_1_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_5_0 <= r_4_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_5_1 <= r_4_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_6_0 <= mesh_1_0_io_out_a_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_6_1 <= mesh_1_0_io_out_a_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_7_0 <= r_6_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_7_1 <= r_6_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    v <= io_in_valid_0_0; // @[Valid.scala 117:22]
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b__0 <= io_in_b_0_0; // @[Reg.scala 16:23]
    end
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b__1 <= io_in_b_0_1; // @[Reg.scala 16:23]
    end
    if (v) begin // @[Reg.scala 16:19]
      outPipe_bits__0 <= b__0; // @[Reg.scala 16:23]
    end
    if (v) begin // @[Reg.scala 16:19]
      outPipe_bits__1 <= b__1; // @[Reg.scala 16:23]
    end
    v_1 <= mesh_0_0_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_1_0 <= mesh_0_0_io_out_b_0; // @[Reg.scala 16:23]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_1_1 <= mesh_0_0_io_out_b_1; // @[Reg.scala 16:23]
    end
    if (v_1) begin // @[Reg.scala 16:19]
      outPipe_bits_1_0 <= b_1_0; // @[Reg.scala 16:23]
    end
    if (v_1) begin // @[Reg.scala 16:19]
      outPipe_bits_1_1 <= b_1_1; // @[Reg.scala 16:23]
    end
    v_2 <= io_in_valid_1_0; // @[Valid.scala 117:22]
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_2_0 <= io_in_b_1_0; // @[Reg.scala 16:23]
    end
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_2_1 <= io_in_b_1_1; // @[Reg.scala 16:23]
    end
    if (v_2) begin // @[Reg.scala 16:19]
      outPipe_bits_2_0 <= b_2_0; // @[Reg.scala 16:23]
    end
    if (v_2) begin // @[Reg.scala 16:19]
      outPipe_bits_2_1 <= b_2_1; // @[Reg.scala 16:23]
    end
    v_3 <= mesh_0_1_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_3_0 <= mesh_0_1_io_out_b_0; // @[Reg.scala 16:23]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_3_1 <= mesh_0_1_io_out_b_1; // @[Reg.scala 16:23]
    end
    if (v_3) begin // @[Reg.scala 16:19]
      outPipe_bits_3_0 <= b_3_0; // @[Reg.scala 16:23]
    end
    if (v_3) begin // @[Reg.scala 16:19]
      outPipe_bits_3_1 <= b_3_1; // @[Reg.scala 16:23]
    end
    v_4 <= io_in_valid_0_0; // @[Valid.scala 117:22]
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b_4_0 <= io_in_d_0_0; // @[Reg.scala 16:23]
    end
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b_4_1 <= io_in_d_0_1; // @[Reg.scala 16:23]
    end
    if (v_4) begin // @[Reg.scala 16:19]
      outPipe_bits_4_0 <= b_4_0; // @[Reg.scala 16:23]
    end
    if (v_4) begin // @[Reg.scala 16:19]
      outPipe_bits_4_1 <= b_4_1; // @[Reg.scala 16:23]
    end
    v_5 <= mesh_0_0_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_5_0 <= mesh_0_0_io_out_c_0; // @[Reg.scala 16:23]
    end
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_5_1 <= mesh_0_0_io_out_c_1; // @[Reg.scala 16:23]
    end
    if (v_5) begin // @[Reg.scala 16:19]
      outPipe_bits_5_0 <= b_5_0; // @[Reg.scala 16:23]
    end
    if (v_5) begin // @[Reg.scala 16:19]
      outPipe_bits_5_1 <= b_5_1; // @[Reg.scala 16:23]
    end
    v_6 <= io_in_valid_1_0; // @[Valid.scala 117:22]
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_6_0 <= io_in_d_1_0; // @[Reg.scala 16:23]
    end
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_6_1 <= io_in_d_1_1; // @[Reg.scala 16:23]
    end
    if (v_6) begin // @[Reg.scala 16:19]
      outPipe_bits_6_0 <= b_6_0; // @[Reg.scala 16:23]
    end
    if (v_6) begin // @[Reg.scala 16:19]
      outPipe_bits_6_1 <= b_6_1; // @[Reg.scala 16:23]
    end
    v_7 <= mesh_0_1_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_7_0 <= mesh_0_1_io_out_c_0; // @[Reg.scala 16:23]
    end
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_7_1 <= mesh_0_1_io_out_c_1; // @[Reg.scala 16:23]
    end
    if (v_7) begin // @[Reg.scala 16:19]
      outPipe_bits_7_0 <= b_7_0; // @[Reg.scala 16:23]
    end
    if (v_7) begin // @[Reg.scala 16:19]
      outPipe_bits_7_1 <= b_7_1; // @[Reg.scala 16:23]
    end
    v_8 <= io_in_valid_0_0; // @[Valid.scala 117:22]
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b_8 <= io_in_control_0_0_shift; // @[Reg.scala 16:23]
    end
    if (v_8) begin // @[Reg.scala 16:19]
      outPipe_bits_8 <= b_8; // @[Reg.scala 16:23]
    end
    v_9 <= io_in_valid_0_0; // @[Valid.scala 117:22]
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b_9 <= io_in_control_0_0_dataflow; // @[Reg.scala 16:23]
    end
    if (v_9) begin // @[Reg.scala 16:19]
      outPipe_bits_9 <= b_9; // @[Reg.scala 16:23]
    end
    v_10 <= io_in_valid_0_0; // @[Valid.scala 117:22]
    if (io_in_valid_0_0) begin // @[Reg.scala 16:19]
      b_10 <= io_in_control_0_0_propagate; // @[Reg.scala 16:23]
    end
    if (v_10) begin // @[Reg.scala 16:19]
      outPipe_bits_10 <= b_10; // @[Reg.scala 16:23]
    end
    v_11 <= io_in_valid_0_1; // @[Valid.scala 117:22]
    if (io_in_valid_0_1) begin // @[Reg.scala 16:19]
      b_11 <= io_in_control_0_1_shift; // @[Reg.scala 16:23]
    end
    if (v_11) begin // @[Reg.scala 16:19]
      outPipe_bits_11 <= b_11; // @[Reg.scala 16:23]
    end
    v_12 <= io_in_valid_0_1; // @[Valid.scala 117:22]
    if (io_in_valid_0_1) begin // @[Reg.scala 16:19]
      b_12 <= io_in_control_0_1_dataflow; // @[Reg.scala 16:23]
    end
    if (v_12) begin // @[Reg.scala 16:19]
      outPipe_bits_12 <= b_12; // @[Reg.scala 16:23]
    end
    v_13 <= io_in_valid_0_1; // @[Valid.scala 117:22]
    if (io_in_valid_0_1) begin // @[Reg.scala 16:19]
      b_13 <= io_in_control_0_1_propagate; // @[Reg.scala 16:23]
    end
    if (v_13) begin // @[Reg.scala 16:19]
      outPipe_bits_13 <= b_13; // @[Reg.scala 16:23]
    end
    v_14 <= mesh_0_0_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_14 <= mesh_0_0_io_out_control_0_shift; // @[Reg.scala 16:23]
    end
    if (v_14) begin // @[Reg.scala 16:19]
      outPipe_bits_14 <= b_14; // @[Reg.scala 16:23]
    end
    v_15 <= mesh_0_0_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_15 <= mesh_0_0_io_out_control_0_dataflow; // @[Reg.scala 16:23]
    end
    if (v_15) begin // @[Reg.scala 16:19]
      outPipe_bits_15 <= b_15; // @[Reg.scala 16:23]
    end
    v_16 <= mesh_0_0_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_16 <= mesh_0_0_io_out_control_0_propagate; // @[Reg.scala 16:23]
    end
    if (v_16) begin // @[Reg.scala 16:19]
      outPipe_bits_16 <= b_16; // @[Reg.scala 16:23]
    end
    v_17 <= mesh_0_0_io_out_valid_1; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_1) begin // @[Reg.scala 16:19]
      b_17 <= mesh_0_0_io_out_control_1_shift; // @[Reg.scala 16:23]
    end
    if (v_17) begin // @[Reg.scala 16:19]
      outPipe_bits_17 <= b_17; // @[Reg.scala 16:23]
    end
    v_18 <= mesh_0_0_io_out_valid_1; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_1) begin // @[Reg.scala 16:19]
      b_18 <= mesh_0_0_io_out_control_1_dataflow; // @[Reg.scala 16:23]
    end
    if (v_18) begin // @[Reg.scala 16:19]
      outPipe_bits_18 <= b_18; // @[Reg.scala 16:23]
    end
    v_19 <= mesh_0_0_io_out_valid_1; // @[Valid.scala 117:22]
    if (mesh_0_0_io_out_valid_1) begin // @[Reg.scala 16:19]
      b_19 <= mesh_0_0_io_out_control_1_propagate; // @[Reg.scala 16:23]
    end
    if (v_19) begin // @[Reg.scala 16:19]
      outPipe_bits_19 <= b_19; // @[Reg.scala 16:23]
    end
    v_20 <= io_in_valid_1_0; // @[Valid.scala 117:22]
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_20 <= io_in_control_1_0_shift; // @[Reg.scala 16:23]
    end
    if (v_20) begin // @[Reg.scala 16:19]
      outPipe_bits_20 <= b_20; // @[Reg.scala 16:23]
    end
    v_21 <= io_in_valid_1_0; // @[Valid.scala 117:22]
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_21 <= io_in_control_1_0_dataflow; // @[Reg.scala 16:23]
    end
    if (v_21) begin // @[Reg.scala 16:19]
      outPipe_bits_21 <= b_21; // @[Reg.scala 16:23]
    end
    v_22 <= io_in_valid_1_0; // @[Valid.scala 117:22]
    if (io_in_valid_1_0) begin // @[Reg.scala 16:19]
      b_22 <= io_in_control_1_0_propagate; // @[Reg.scala 16:23]
    end
    if (v_22) begin // @[Reg.scala 16:19]
      outPipe_bits_22 <= b_22; // @[Reg.scala 16:23]
    end
    v_23 <= io_in_valid_1_1; // @[Valid.scala 117:22]
    if (io_in_valid_1_1) begin // @[Reg.scala 16:19]
      b_23 <= io_in_control_1_1_shift; // @[Reg.scala 16:23]
    end
    if (v_23) begin // @[Reg.scala 16:19]
      outPipe_bits_23 <= b_23; // @[Reg.scala 16:23]
    end
    v_24 <= io_in_valid_1_1; // @[Valid.scala 117:22]
    if (io_in_valid_1_1) begin // @[Reg.scala 16:19]
      b_24 <= io_in_control_1_1_dataflow; // @[Reg.scala 16:23]
    end
    if (v_24) begin // @[Reg.scala 16:19]
      outPipe_bits_24 <= b_24; // @[Reg.scala 16:23]
    end
    v_25 <= io_in_valid_1_1; // @[Valid.scala 117:22]
    if (io_in_valid_1_1) begin // @[Reg.scala 16:19]
      b_25 <= io_in_control_1_1_propagate; // @[Reg.scala 16:23]
    end
    if (v_25) begin // @[Reg.scala 16:19]
      outPipe_bits_25 <= b_25; // @[Reg.scala 16:23]
    end
    v_26 <= mesh_0_1_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_26 <= mesh_0_1_io_out_control_0_shift; // @[Reg.scala 16:23]
    end
    if (v_26) begin // @[Reg.scala 16:19]
      outPipe_bits_26 <= b_26; // @[Reg.scala 16:23]
    end
    v_27 <= mesh_0_1_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_27 <= mesh_0_1_io_out_control_0_dataflow; // @[Reg.scala 16:23]
    end
    if (v_27) begin // @[Reg.scala 16:19]
      outPipe_bits_27 <= b_27; // @[Reg.scala 16:23]
    end
    v_28 <= mesh_0_1_io_out_valid_0; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_0) begin // @[Reg.scala 16:19]
      b_28 <= mesh_0_1_io_out_control_0_propagate; // @[Reg.scala 16:23]
    end
    if (v_28) begin // @[Reg.scala 16:19]
      outPipe_bits_28 <= b_28; // @[Reg.scala 16:23]
    end
    v_29 <= mesh_0_1_io_out_valid_1; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_1) begin // @[Reg.scala 16:19]
      b_29 <= mesh_0_1_io_out_control_1_shift; // @[Reg.scala 16:23]
    end
    if (v_29) begin // @[Reg.scala 16:19]
      outPipe_bits_29 <= b_29; // @[Reg.scala 16:23]
    end
    v_30 <= mesh_0_1_io_out_valid_1; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_1) begin // @[Reg.scala 16:19]
      b_30 <= mesh_0_1_io_out_control_1_dataflow; // @[Reg.scala 16:23]
    end
    if (v_30) begin // @[Reg.scala 16:19]
      outPipe_bits_30 <= b_30; // @[Reg.scala 16:23]
    end
    v_31 <= mesh_0_1_io_out_valid_1; // @[Valid.scala 117:22]
    if (mesh_0_1_io_out_valid_1) begin // @[Reg.scala 16:19]
      b_31 <= mesh_0_1_io_out_control_1_propagate; // @[Reg.scala 16:23]
    end
    if (v_31) begin // @[Reg.scala 16:19]
      outPipe_bits_31 <= b_31; // @[Reg.scala 16:23]
    end
    r_8_0 <= io_in_valid_0_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_8_1 <= io_in_valid_0_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_9_0 <= r_8_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_9_1 <= r_8_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_10_0 <= mesh_0_0_io_out_valid_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_10_1 <= mesh_0_0_io_out_valid_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_11_0 <= r_10_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_11_1 <= r_10_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_12_0 <= io_in_valid_1_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_12_1 <= io_in_valid_1_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_13_0 <= r_12_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_13_1 <= r_12_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_14_0 <= mesh_0_1_io_out_valid_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_14_1 <= mesh_0_1_io_out_valid_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_15_0 <= r_14_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_15_1 <= r_14_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_16_0 <= io_in_id_0_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_16_1 <= io_in_id_0_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_17_0 <= r_16_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_17_1 <= r_16_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_18_0 <= mesh_0_0_io_out_id_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_18_1 <= mesh_0_0_io_out_id_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_19_0 <= r_18_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_19_1 <= r_18_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_20_0 <= io_in_id_1_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_20_1 <= io_in_id_1_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_21_0 <= r_20_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_21_1 <= r_20_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_22_0 <= mesh_0_1_io_out_id_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_22_1 <= mesh_0_1_io_out_id_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_23_0 <= r_22_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_23_1 <= r_22_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_24_0 <= io_in_last_0_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_24_1 <= io_in_last_0_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_25_0 <= r_24_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_25_1 <= r_24_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_26_0 <= mesh_0_0_io_out_last_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_26_1 <= mesh_0_0_io_out_last_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_27_0 <= r_26_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_27_1 <= r_26_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_28_0 <= io_in_last_1_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_28_1 <= io_in_last_1_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_29_0 <= r_28_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_29_1 <= r_28_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_30_0 <= mesh_0_1_io_out_last_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_30_1 <= mesh_0_1_io_out_last_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_31_0 <= r_30_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_31_1 <= r_30_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_32_0 <= mesh_1_0_io_out_b_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_32_1 <= mesh_1_0_io_out_b_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_33_0 <= mesh_1_0_io_out_c_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_33_1 <= mesh_1_0_io_out_c_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_34_0 <= mesh_1_0_io_out_valid_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_35_0_dataflow <= mesh_1_0_io_out_control_0_dataflow; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_36_0 <= mesh_1_0_io_out_id_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_37_0 <= mesh_1_0_io_out_last_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_38_0 <= mesh_1_1_io_out_b_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_38_1 <= mesh_1_1_io_out_b_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_39_0 <= mesh_1_1_io_out_c_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_39_1 <= mesh_1_1_io_out_c_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r__0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  r__1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  r_1_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  r_1_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  r_2_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  r_2_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  r_3_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  r_3_1 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  r_4_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  r_4_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  r_5_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  r_5_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  r_6_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  r_6_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  r_7_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  r_7_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  v = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  b__0 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  b__1 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  outPipe_bits__0 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  outPipe_bits__1 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  v_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  b_1_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  b_1_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  outPipe_bits_1_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  outPipe_bits_1_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  v_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  b_2_0 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  b_2_1 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  outPipe_bits_2_0 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  outPipe_bits_2_1 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  v_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  b_3_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  b_3_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  outPipe_bits_3_0 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  outPipe_bits_3_1 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  v_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  b_4_0 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  b_4_1 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  outPipe_bits_4_0 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  outPipe_bits_4_1 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  v_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  b_5_0 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  b_5_1 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  outPipe_bits_5_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  outPipe_bits_5_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  v_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  b_6_0 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  b_6_1 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  outPipe_bits_6_0 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  outPipe_bits_6_1 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  v_7 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  b_7_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  b_7_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  outPipe_bits_7_0 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  outPipe_bits_7_1 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  v_8 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  b_8 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  outPipe_bits_8 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  v_9 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  b_9 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  outPipe_bits_9 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  v_10 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  b_10 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  outPipe_bits_10 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  v_11 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  b_11 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  outPipe_bits_11 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  v_12 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  b_12 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  outPipe_bits_12 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  v_13 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  b_13 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  outPipe_bits_13 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  v_14 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  b_14 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  outPipe_bits_14 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  v_15 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  b_15 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  outPipe_bits_15 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  v_16 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  b_16 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  outPipe_bits_16 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  v_17 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  b_17 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  outPipe_bits_17 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  v_18 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  b_18 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  outPipe_bits_18 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  v_19 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  b_19 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  outPipe_bits_19 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  v_20 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  b_20 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  outPipe_bits_20 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  v_21 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  b_21 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  outPipe_bits_21 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  v_22 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  b_22 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  outPipe_bits_22 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  v_23 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  b_23 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  outPipe_bits_23 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  v_24 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  b_24 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  outPipe_bits_24 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  v_25 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  b_25 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  outPipe_bits_25 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  v_26 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  b_26 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  outPipe_bits_26 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  v_27 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  b_27 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  outPipe_bits_27 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  v_28 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  b_28 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  outPipe_bits_28 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  v_29 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  b_29 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  outPipe_bits_29 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  v_30 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  b_30 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  outPipe_bits_30 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  v_31 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  b_31 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  outPipe_bits_31 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r_8_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r_8_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r_9_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r_9_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r_10_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r_10_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r_11_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r_11_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r_12_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r_12_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_13_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_13_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_14_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_14_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_15_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_15_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_16_0 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  r_16_1 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  r_17_0 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  r_17_1 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  r_18_0 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  r_18_1 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  r_19_0 = _RAND_150[2:0];
  _RAND_151 = {1{`RANDOM}};
  r_19_1 = _RAND_151[2:0];
  _RAND_152 = {1{`RANDOM}};
  r_20_0 = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  r_20_1 = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  r_21_0 = _RAND_154[2:0];
  _RAND_155 = {1{`RANDOM}};
  r_21_1 = _RAND_155[2:0];
  _RAND_156 = {1{`RANDOM}};
  r_22_0 = _RAND_156[2:0];
  _RAND_157 = {1{`RANDOM}};
  r_22_1 = _RAND_157[2:0];
  _RAND_158 = {1{`RANDOM}};
  r_23_0 = _RAND_158[2:0];
  _RAND_159 = {1{`RANDOM}};
  r_23_1 = _RAND_159[2:0];
  _RAND_160 = {1{`RANDOM}};
  r_24_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_24_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_25_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_25_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_26_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_26_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_27_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r_27_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r_28_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r_28_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r_29_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r_29_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r_30_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r_30_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r_31_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r_31_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r_32_0 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  r_32_1 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  r_33_0 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  r_33_1 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  r_34_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r_35_0_dataflow = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r_36_0 = _RAND_182[2:0];
  _RAND_183 = {1{`RANDOM}};
  r_37_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r_38_0 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  r_38_1 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  r_39_0 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  r_39_1 = _RAND_187[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TagQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_tag,
  input  [2:0]  io_enq_bits_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_tag,
  output [2:0]  io_deq_bits_id,
  output [31:0] io_all_0_tag,
  output [31:0] io_all_1_tag,
  output [31:0] io_all_2_tag,
  output [31:0] io_all_3_tag,
  output [31:0] io_all_4_tag,
  output [31:0] io_all_5_tag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0_tag; // @[TagQueue.scala 18:17]
  reg [2:0] regs_0_id; // @[TagQueue.scala 18:17]
  reg [31:0] regs_1_tag; // @[TagQueue.scala 18:17]
  reg [2:0] regs_1_id; // @[TagQueue.scala 18:17]
  reg [31:0] regs_2_tag; // @[TagQueue.scala 18:17]
  reg [2:0] regs_2_id; // @[TagQueue.scala 18:17]
  reg [31:0] regs_3_tag; // @[TagQueue.scala 18:17]
  reg [2:0] regs_3_id; // @[TagQueue.scala 18:17]
  reg [31:0] regs_4_tag; // @[TagQueue.scala 18:17]
  reg [2:0] regs_4_id; // @[TagQueue.scala 18:17]
  reg [31:0] regs_5_tag; // @[TagQueue.scala 18:17]
  reg [2:0] regs_5_id; // @[TagQueue.scala 18:17]
  reg [2:0] raddr; // @[TagQueue.scala 19:22]
  reg [2:0] waddr; // @[TagQueue.scala 20:22]
  reg [2:0] len; // @[TagQueue.scala 21:20]
  wire  empty = len == 3'h0; // @[TagQueue.scala 23:19]
  wire  full = len == 3'h6; // @[TagQueue.scala 24:18]
  wire [2:0] _GEN_7 = 3'h1 == raddr ? regs_1_id : regs_0_id; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [2:0] _GEN_8 = 3'h2 == raddr ? regs_2_id : _GEN_7; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [2:0] _GEN_9 = 3'h3 == raddr ? regs_3_id : _GEN_8; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [2:0] _GEN_10 = 3'h4 == raddr ? regs_4_id : _GEN_9; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [31:0] _GEN_13 = 3'h1 == raddr ? regs_1_tag : regs_0_tag; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [31:0] _GEN_14 = 3'h2 == raddr ? regs_2_tag : _GEN_13; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [31:0] _GEN_15 = 3'h3 == raddr ? regs_3_tag : _GEN_14; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire [31:0] _GEN_16 = 3'h4 == raddr ? regs_4_tag : _GEN_15; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  wire  _T_2 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_8 = 3'h5 - 3'h1; // @[Util.scala 13:22]
  wire [2:0] _T_10 = _T_8 + 3'h1; // @[Util.scala 13:26]
  wire [2:0] _T_15 = 3'h5 - waddr; // @[Util.scala 13:57]
  wire [2:0] _T_17 = 3'h1 - _T_15; // @[Util.scala 13:48]
  wire [2:0] _T_19 = _T_17 - 3'h1; // @[Util.scala 13:62]
  wire [2:0] _T_21 = waddr + 3'h1; // @[Util.scala 13:71]
  wire  _T_23 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_36 = 3'h5 - raddr; // @[Util.scala 13:57]
  wire [2:0] _T_38 = 3'h1 - _T_36; // @[Util.scala 13:48]
  wire [2:0] _T_40 = _T_38 - 3'h1; // @[Util.scala 13:62]
  wire [2:0] _T_42 = raddr + 3'h1; // @[Util.scala 13:71]
  wire [2:0] _T_49 = len + 3'h1; // @[TagQueue.scala 42:16]
  wire [2:0] _T_55 = len - 3'h1; // @[TagQueue.scala 44:16]
  assign io_enq_ready = ~full; // @[TagQueue.scala 26:19]
  assign io_deq_valid = ~empty; // @[TagQueue.scala 27:19]
  assign io_deq_bits_tag = 3'h5 == raddr ? regs_5_tag : _GEN_16; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  assign io_deq_bits_id = 3'h5 == raddr ? regs_5_id : _GEN_10; // @[TagQueue.scala 28:15 TagQueue.scala 28:15]
  assign io_all_0_tag = regs_0_tag; // @[TagQueue.scala 29:10]
  assign io_all_1_tag = regs_1_tag; // @[TagQueue.scala 29:10]
  assign io_all_2_tag = regs_2_tag; // @[TagQueue.scala 29:10]
  assign io_all_3_tag = regs_3_tag; // @[TagQueue.scala 29:10]
  assign io_all_4_tag = regs_4_tag; // @[TagQueue.scala 29:10]
  assign io_all_5_tag = regs_5_tag; // @[TagQueue.scala 29:10]
  always @(posedge clock) begin
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h0 == waddr) begin // @[TagQueue.scala 32:17]
        regs_0_tag <= io_enq_bits_tag; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h0 == waddr) begin // @[TagQueue.scala 32:17]
        regs_0_id <= io_enq_bits_id; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h1 == waddr) begin // @[TagQueue.scala 32:17]
        regs_1_tag <= io_enq_bits_tag; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h1 == waddr) begin // @[TagQueue.scala 32:17]
        regs_1_id <= io_enq_bits_id; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h2 == waddr) begin // @[TagQueue.scala 32:17]
        regs_2_tag <= io_enq_bits_tag; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h2 == waddr) begin // @[TagQueue.scala 32:17]
        regs_2_id <= io_enq_bits_id; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h3 == waddr) begin // @[TagQueue.scala 32:17]
        regs_3_tag <= io_enq_bits_tag; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h3 == waddr) begin // @[TagQueue.scala 32:17]
        regs_3_id <= io_enq_bits_id; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h4 == waddr) begin // @[TagQueue.scala 32:17]
        regs_4_tag <= io_enq_bits_tag; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h4 == waddr) begin // @[TagQueue.scala 32:17]
        regs_4_id <= io_enq_bits_id; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h5 == waddr) begin // @[TagQueue.scala 32:17]
        regs_5_tag <= io_enq_bits_tag; // @[TagQueue.scala 32:17]
      end
    end
    if (_T_2) begin // @[TagQueue.scala 31:22]
      if (3'h5 == waddr) begin // @[TagQueue.scala 32:17]
        regs_5_id <= io_enq_bits_id; // @[TagQueue.scala 32:17]
      end
    end
    if (reset) begin // @[TagQueue.scala 19:22]
      raddr <= 3'h0; // @[TagQueue.scala 19:22]
    end else if (_T_23) begin // @[TagQueue.scala 36:22]
      if (raddr >= _T_10) begin // @[Util.scala 13:10]
        raddr <= _T_40;
      end else begin
        raddr <= _T_42;
      end
    end
    if (reset) begin // @[TagQueue.scala 20:22]
      waddr <= 3'h0; // @[TagQueue.scala 20:22]
    end else if (_T_2) begin // @[TagQueue.scala 31:22]
      if (waddr >= _T_10) begin // @[Util.scala 13:10]
        waddr <= _T_19;
      end else begin
        waddr <= _T_21;
      end
    end
    if (reset) begin // @[TagQueue.scala 21:20]
      len <= 3'h0; // @[TagQueue.scala 21:20]
    end else if (_T_2 & ~_T_23) begin // @[TagQueue.scala 41:38]
      len <= _T_49; // @[TagQueue.scala 42:9]
    end else if (~_T_2 & _T_23) begin // @[TagQueue.scala 43:43]
      len <= _T_55; // @[TagQueue.scala 44:9]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(len <= 3'h6 | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TagQueue.scala:51 assert(len <= entries.U)\n"); // @[TagQueue.scala 51:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(len <= 3'h6 | reset)) begin
          $fatal; // @[TagQueue.scala 51:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0_tag = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_0_id = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  regs_1_tag = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_1_id = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  regs_2_tag = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_2_id = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  regs_3_tag = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_3_id = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  regs_4_tag = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_4_id = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  regs_5_tag = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_5_id = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  raddr = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  waddr = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  len = _RAND_14[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_id,
  input  [2:0] io_enq_bits_total_rows,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_id,
  output [2:0] io_deq_bits_total_rows
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] ram_id [0:5]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_total_rows [0:5]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_total_rows_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_total_rows_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_total_rows_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_total_rows_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_total_rows_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_total_rows_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 3'h5; // @[Counter.scala 72:24]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  wire  wrap_1 = deq_ptr_value == 3'h5; // @[Counter.scala 72:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  assign ram_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_id_io_deq_bits_MPORT_data = ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_id_io_deq_bits_MPORT_data = ram_id_io_deq_bits_MPORT_addr >= 3'h6 ? _RAND_1[2:0] :
    ram_id[ram_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_id_MPORT_data = io_enq_bits_id;
  assign ram_id_MPORT_addr = enq_ptr_value;
  assign ram_id_MPORT_mask = 1'h1;
  assign ram_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_total_rows_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_total_rows_io_deq_bits_MPORT_data = ram_total_rows[ram_total_rows_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_total_rows_io_deq_bits_MPORT_data = ram_total_rows_io_deq_bits_MPORT_addr >= 3'h6 ? _RAND_3[2:0] :
    ram_total_rows[ram_total_rows_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_total_rows_MPORT_data = io_enq_bits_total_rows;
  assign ram_total_rows_MPORT_addr = enq_ptr_value;
  assign ram_total_rows_MPORT_mask = 1'h1;
  assign ram_total_rows_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_id = ram_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_total_rows = ram_total_rows_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_id_MPORT_en & ram_id_MPORT_mask) begin
      ram_id[ram_id_MPORT_addr] <= ram_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_total_rows_MPORT_en & ram_total_rows_MPORT_mask) begin
      ram_total_rows[ram_total_rows_MPORT_addr] <= ram_total_rows_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      if (wrap) begin // @[Counter.scala 86:20]
        enq_ptr_value <= 3'h0; // @[Counter.scala 86:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      if (wrap_1) begin // @[Counter.scala 86:20]
        deq_ptr_value <= 3'h0; // @[Counter.scala 86:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[2:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    ram_total_rows[initvar] = _RAND_2[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enq_ptr_value = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  deq_ptr_value = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  maybe_full = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MeshWithDelays(
  input         clock,
  input         reset,
  output        io_a_ready,
  input         io_a_valid,
  input  [7:0]  io_a_bits_0_0,
  input  [7:0]  io_a_bits_0_1,
  input  [7:0]  io_a_bits_1_0,
  input  [7:0]  io_a_bits_1_1,
  output        io_b_ready,
  input         io_b_valid,
  input  [7:0]  io_b_bits_0_0,
  input  [7:0]  io_b_bits_0_1,
  input  [7:0]  io_b_bits_1_0,
  input  [7:0]  io_b_bits_1_1,
  output        io_d_ready,
  input         io_d_valid,
  input  [7:0]  io_d_bits_0_0,
  input  [7:0]  io_d_bits_0_1,
  input  [7:0]  io_d_bits_1_0,
  input  [7:0]  io_d_bits_1_1,
  output        io_req_ready,
  input         io_req_valid,
  input         io_req_bits_pe_control_dataflow,
  input         io_req_bits_pe_control_propagate,
  input  [3:0]  io_req_bits_pe_control_shift,
  input         io_req_bits_a_transpose,
  input         io_req_bits_bd_transpose,
  input  [2:0]  io_req_bits_total_rows,
  input  [31:0] io_req_bits_tag,
  input  [1:0]  io_req_bits_flush,
  output        io_resp_valid,
  output [7:0]  io_resp_bits_data_0_0,
  output [7:0]  io_resp_bits_data_0_1,
  output [7:0]  io_resp_bits_data_1_0,
  output [7:0]  io_resp_bits_data_1_1,
  output [2:0]  io_resp_bits_total_rows,
  output [31:0] io_resp_bits_tag,
  output        io_resp_bits_last,
  output [31:0] io_tags_in_progress_0,
  output [31:0] io_tags_in_progress_1,
  output [31:0] io_tags_in_progress_2,
  output [31:0] io_tags_in_progress_3,
  output [31:0] io_tags_in_progress_4,
  output [31:0] io_tags_in_progress_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
`endif // RANDOMIZE_REG_INIT
  wire  transposer_clock; // @[MeshWithDelays.scala 154:26]
  wire  transposer_reset; // @[MeshWithDelays.scala 154:26]
  wire  transposer_io_inRow_ready; // @[MeshWithDelays.scala 154:26]
  wire  transposer_io_inRow_valid; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_inRow_bits_0; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_inRow_bits_1; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_inRow_bits_2; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_inRow_bits_3; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_outCol_bits_0; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_outCol_bits_1; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_outCol_bits_2; // @[MeshWithDelays.scala 154:26]
  wire [7:0] transposer_io_outCol_bits_3; // @[MeshWithDelays.scala 154:26]
  wire  mesh_clock; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_a_0_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_a_0_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_a_1_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_a_1_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_b_0_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_b_0_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_b_1_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_b_1_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_d_0_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_d_0_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_d_1_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_in_d_1_1; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_0_0_dataflow; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_0_0_propagate; // @[MeshWithDelays.scala 166:20]
  wire [3:0] mesh_io_in_control_0_0_shift; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_0_1_dataflow; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_0_1_propagate; // @[MeshWithDelays.scala 166:20]
  wire [3:0] mesh_io_in_control_0_1_shift; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_1_0_dataflow; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_1_0_propagate; // @[MeshWithDelays.scala 166:20]
  wire [3:0] mesh_io_in_control_1_0_shift; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_1_1_dataflow; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_control_1_1_propagate; // @[MeshWithDelays.scala 166:20]
  wire [3:0] mesh_io_in_control_1_1_shift; // @[MeshWithDelays.scala 166:20]
  wire [2:0] mesh_io_in_id_0_0; // @[MeshWithDelays.scala 166:20]
  wire [2:0] mesh_io_in_id_0_1; // @[MeshWithDelays.scala 166:20]
  wire [2:0] mesh_io_in_id_1_0; // @[MeshWithDelays.scala 166:20]
  wire [2:0] mesh_io_in_id_1_1; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_last_0_0; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_last_0_1; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_last_1_0; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_last_1_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_b_0_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_b_0_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_b_1_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_b_1_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_c_0_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_c_0_1; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_c_1_0; // @[MeshWithDelays.scala 166:20]
  wire [7:0] mesh_io_out_c_1_1; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_valid_0_0; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_valid_0_1; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_valid_1_0; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_in_valid_1_1; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_out_valid_0_0; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_out_control_0_0_dataflow; // @[MeshWithDelays.scala 166:20]
  wire [2:0] mesh_io_out_id_0_0; // @[MeshWithDelays.scala 166:20]
  wire  mesh_io_out_last_0_0; // @[MeshWithDelays.scala 166:20]
  wire  tagq_clock; // @[MeshWithDelays.scala 221:20]
  wire  tagq_reset; // @[MeshWithDelays.scala 221:20]
  wire  tagq_io_enq_ready; // @[MeshWithDelays.scala 221:20]
  wire  tagq_io_enq_valid; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_enq_bits_tag; // @[MeshWithDelays.scala 221:20]
  wire [2:0] tagq_io_enq_bits_id; // @[MeshWithDelays.scala 221:20]
  wire  tagq_io_deq_ready; // @[MeshWithDelays.scala 221:20]
  wire  tagq_io_deq_valid; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_deq_bits_tag; // @[MeshWithDelays.scala 221:20]
  wire [2:0] tagq_io_deq_bits_id; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_all_0_tag; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_all_1_tag; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_all_2_tag; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_all_3_tag; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_all_4_tag; // @[MeshWithDelays.scala 221:20]
  wire [31:0] tagq_io_all_5_tag; // @[MeshWithDelays.scala 221:20]
  wire  total_rows_q_clock; // @[MeshWithDelays.scala 238:28]
  wire  total_rows_q_reset; // @[MeshWithDelays.scala 238:28]
  wire  total_rows_q_io_enq_ready; // @[MeshWithDelays.scala 238:28]
  wire  total_rows_q_io_enq_valid; // @[MeshWithDelays.scala 238:28]
  wire [2:0] total_rows_q_io_enq_bits_id; // @[MeshWithDelays.scala 238:28]
  wire [2:0] total_rows_q_io_enq_bits_total_rows; // @[MeshWithDelays.scala 238:28]
  wire  total_rows_q_io_deq_ready; // @[MeshWithDelays.scala 238:28]
  wire  total_rows_q_io_deq_valid; // @[MeshWithDelays.scala 238:28]
  wire [2:0] total_rows_q_io_deq_bits_id; // @[MeshWithDelays.scala 238:28]
  wire [2:0] total_rows_q_io_deq_bits_total_rows; // @[MeshWithDelays.scala 238:28]
  reg  req_valid; // @[MeshWithDelays.scala 92:16]
  reg  req_bits_pe_control_dataflow; // @[MeshWithDelays.scala 92:16]
  reg [3:0] req_bits_pe_control_shift; // @[MeshWithDelays.scala 92:16]
  reg  req_bits_a_transpose; // @[MeshWithDelays.scala 92:16]
  reg  req_bits_bd_transpose; // @[MeshWithDelays.scala 92:16]
  reg [2:0] req_bits_total_rows; // @[MeshWithDelays.scala 92:16]
  reg [1:0] req_bits_flush; // @[MeshWithDelays.scala 92:16]
  reg [2:0] matmul_id; // @[MeshWithDelays.scala 94:26]
  reg [1:0] fire_counter; // @[MeshWithDelays.scala 97:29]
  wire  _T = io_a_ready & io_a_valid; // @[Decoupled.scala 40:37]
  reg [7:0] a_buf_0_0; // @[Reg.scala 15:16]
  reg [7:0] a_buf_0_1; // @[Reg.scala 15:16]
  reg [7:0] a_buf_1_0; // @[Reg.scala 15:16]
  reg [7:0] a_buf_1_1; // @[Reg.scala 15:16]
  wire  _T_1 = io_b_ready & io_b_valid; // @[Decoupled.scala 40:37]
  reg [7:0] b_buf_0_0; // @[Reg.scala 15:16]
  reg [7:0] b_buf_0_1; // @[Reg.scala 15:16]
  reg [7:0] b_buf_1_0; // @[Reg.scala 15:16]
  reg [7:0] b_buf_1_1; // @[Reg.scala 15:16]
  wire  _T_2 = io_d_ready & io_d_valid; // @[Decoupled.scala 40:37]
  reg [7:0] d_buf_0_0; // @[Reg.scala 15:16]
  reg [7:0] d_buf_0_1; // @[Reg.scala 15:16]
  reg [7:0] d_buf_1_0; // @[Reg.scala 15:16]
  reg [7:0] d_buf_1_1; // @[Reg.scala 15:16]
  reg  a_written; // @[MeshWithDelays.scala 103:26]
  reg  b_written; // @[MeshWithDelays.scala 104:26]
  reg  d_written; // @[MeshWithDelays.scala 105:26]
  reg  in_prop; // @[MeshWithDelays.scala 107:20]
  wire  input_next_row_into_spatial_array = req_valid & (a_written & b_written & d_written | req_bits_flush > 2'h0); // @[MeshWithDelays.scala 109:53]
  wire [2:0] _T_8 = req_bits_total_rows - 3'h1; // @[MeshWithDelays.scala 111:48]
  wire [2:0] _GEN_85 = {{1'd0}, fire_counter}; // @[MeshWithDelays.scala 111:32]
  wire  last_fire = _GEN_85 == _T_8 & input_next_row_into_spatial_array; // @[MeshWithDelays.scala 111:54]
  wire  _T_10 = io_req_ready & io_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_17 = 3'h4 - 3'h1; // @[Util.scala 13:22]
  wire [2:0] _T_19 = _T_17 + 3'h1; // @[Util.scala 13:26]
  wire [2:0] _T_24 = 3'h4 - matmul_id; // @[Util.scala 13:57]
  wire [2:0] _T_26 = 3'h1 - _T_24; // @[Util.scala 13:48]
  wire [2:0] _T_28 = _T_26 - 3'h1; // @[Util.scala 13:62]
  wire [2:0] _T_30 = matmul_id + 3'h1; // @[Util.scala 13:71]
  wire [1:0] _T_34 = req_bits_flush - 2'h1; // @[MeshWithDelays.scala 119:38]
  wire  _GEN_12 = last_fire ? req_bits_flush > 2'h1 : req_valid; // @[MeshWithDelays.scala 117:26 MeshWithDelays.scala 118:15 MeshWithDelays.scala 92:16]
  wire  _GEN_14 = _T_10 | _GEN_12; // @[MeshWithDelays.scala 113:22 Util.scala 134:13]
  wire  _T_38 = _T_8 == 3'h0; // @[Util.scala 19:28]
  wire [1:0] _T_44 = fire_counter + 2'h1; // @[Util.scala 27:15]
  wire [2:0] _T_48 = _T_8 - 3'h1; // @[Util.scala 30:17]
  wire [2:0] _T_50 = _T_48 + 3'h1; // @[Util.scala 30:21]
  wire  _T_51 = _GEN_85 >= _T_50; // @[Util.scala 30:10]
  wire [2:0] _T_55 = _T_8 - _GEN_85; // @[Util.scala 30:54]
  wire [2:0] _T_57 = 3'h1 - _T_55; // @[Util.scala 30:47]
  wire [2:0] _T_59 = _T_57 - 3'h1; // @[Util.scala 30:59]
  wire [2:0] _T_60 = _T_51 ? _T_59 : {{1'd0}, _T_44}; // @[Mux.scala 98:16]
  wire [2:0] _T_61 = _T_38 ? 3'h0 : _T_60; // @[Mux.scala 98:16]
  wire  _GEN_25 = input_next_row_into_spatial_array ? 1'h0 : a_written; // @[MeshWithDelays.scala 122:44 MeshWithDelays.scala 123:15 MeshWithDelays.scala 103:26]
  wire  _GEN_26 = input_next_row_into_spatial_array ? 1'h0 : b_written; // @[MeshWithDelays.scala 122:44 MeshWithDelays.scala 124:15 MeshWithDelays.scala 104:26]
  wire  _GEN_27 = input_next_row_into_spatial_array ? 1'h0 : d_written; // @[MeshWithDelays.scala 122:44 MeshWithDelays.scala 125:15 MeshWithDelays.scala 105:26]
  wire [2:0] _GEN_28 = input_next_row_into_spatial_array ? _T_61 : {{1'd0}, fire_counter}; // @[MeshWithDelays.scala 122:44 MeshWithDelays.scala 127:18 MeshWithDelays.scala 97:29]
  wire  _GEN_29 = _T | _GEN_25; // @[MeshWithDelays.scala 130:20 MeshWithDelays.scala 131:15]
  wire  _GEN_30 = _T_1 | _GEN_26; // @[MeshWithDelays.scala 134:20 MeshWithDelays.scala 135:15]
  wire  _GEN_31 = _T_2 | _GEN_27; // @[MeshWithDelays.scala 138:20 MeshWithDelays.scala 139:15]
  wire  _T_75 = ~input_next_row_into_spatial_array; // @[MeshWithDelays.scala 146:23]
  wire  _T_80 = ~req_valid; // @[MeshWithDelays.scala 148:15]
  wire  pause = ~req_valid | _T_75; // @[MeshWithDelays.scala 148:26]
  wire  _T_82 = ~req_bits_pe_control_dataflow; // @[MeshWithDelays.scala 151:63]
  wire  a_is_from_transposer = ~req_bits_pe_control_dataflow ? ~req_bits_a_transpose : req_bits_a_transpose; // @[MeshWithDelays.scala 151:33]
  wire  b_is_from_transposer = _T_82 & req_bits_bd_transpose; // @[MeshWithDelays.scala 152:80]
  wire  d_is_from_transposer = req_bits_pe_control_dataflow & req_bits_bd_transpose; // @[MeshWithDelays.scala 153:80]
  wire [7:0] _T_90_0 = d_is_from_transposer ? $signed(d_buf_1_1) : $signed(a_buf_0_0); // @[Mux.scala 98:16]
  wire [7:0] _T_90_1 = d_is_from_transposer ? $signed(d_buf_1_0) : $signed(a_buf_0_1); // @[Mux.scala 98:16]
  wire [7:0] _T_90_2 = d_is_from_transposer ? $signed(d_buf_0_1) : $signed(a_buf_1_0); // @[Mux.scala 98:16]
  wire [7:0] _T_90_3 = d_is_from_transposer ? $signed(d_buf_0_0) : $signed(a_buf_1_1); // @[Mux.scala 98:16]
  wire [31:0] _T_96 = {transposer_io_outCol_bits_3,transposer_io_outCol_bits_2,transposer_io_outCol_bits_1,
    transposer_io_outCol_bits_0}; // @[MeshWithDelays.scala 169:80]
  wire [7:0] _T_98 = _T_96[7:0]; // @[MeshWithDelays.scala 169:80]
  wire [7:0] _T_100 = _T_96[15:8]; // @[MeshWithDelays.scala 169:80]
  wire [7:0] _T_102 = _T_96[23:16]; // @[MeshWithDelays.scala 169:80]
  wire [7:0] _T_104 = _T_96[31:24]; // @[MeshWithDelays.scala 169:80]
  wire [31:0] _T_124 = {transposer_io_outCol_bits_0,transposer_io_outCol_bits_1,transposer_io_outCol_bits_2,
    transposer_io_outCol_bits_3}; // @[MeshWithDelays.scala 172:93]
  wire [7:0] _T_126 = _T_124[7:0]; // @[MeshWithDelays.scala 172:93]
  wire [7:0] _T_128 = _T_124[15:8]; // @[MeshWithDelays.scala 172:93]
  wire [7:0] _T_130 = _T_124[23:16]; // @[MeshWithDelays.scala 172:93]
  wire [7:0] _T_132 = _T_124[31:24]; // @[MeshWithDelays.scala 172:93]
  reg [7:0] r__0; // @[Reg.scala 15:16]
  reg [7:0] r__1; // @[Reg.scala 15:16]
  reg [7:0] r_1_0; // @[Reg.scala 15:16]
  reg [7:0] r_1_1; // @[Reg.scala 15:16]
  reg [7:0] r_2_0; // @[Reg.scala 15:16]
  reg [7:0] r_2_1; // @[Reg.scala 15:16]
  reg [7:0] r_3_0; // @[Reg.scala 15:16]
  reg [7:0] r_3_1; // @[Reg.scala 15:16]
  reg [7:0] r_4_0; // @[Reg.scala 15:16]
  reg [7:0] r_4_1; // @[Reg.scala 15:16]
  reg [7:0] r_5_0; // @[Reg.scala 15:16]
  reg [7:0] r_5_1; // @[Reg.scala 15:16]
  reg  r_6; // @[Reg.scala 15:16]
  reg  r_7; // @[Reg.scala 15:16]
  reg  r_8; // @[Reg.scala 15:16]
  reg  r_9; // @[Reg.scala 15:16]
  reg  r_10; // @[Reg.scala 15:16]
  reg  r_11; // @[Reg.scala 15:16]
  reg  r_12; // @[Reg.scala 15:16]
  reg  r_13; // @[Reg.scala 15:16]
  reg [3:0] result_shift; // @[MeshWithDelays.scala 182:29]
  reg [3:0] r_14; // @[Reg.scala 15:16]
  reg [3:0] r_15; // @[Reg.scala 15:16]
  reg [3:0] r_16; // @[Reg.scala 15:16]
  reg [3:0] r_17; // @[Reg.scala 15:16]
  reg  r_18_0; // @[Reg.scala 15:16]
  reg  r_18_1; // @[Reg.scala 15:16]
  reg  r_19_0; // @[Reg.scala 15:16]
  reg  r_19_1; // @[Reg.scala 15:16]
  reg [2:0] r_20_0; // @[Reg.scala 15:16]
  reg [2:0] r_20_1; // @[Reg.scala 15:16]
  reg [2:0] r_21_0; // @[Reg.scala 15:16]
  reg [2:0] r_21_1; // @[Reg.scala 15:16]
  reg  r_22_0; // @[Reg.scala 15:16]
  reg  r_22_1; // @[Reg.scala 15:16]
  reg  r_23_0; // @[Reg.scala 15:16]
  reg  r_23_1; // @[Reg.scala 15:16]
  reg [7:0] r_24_0; // @[Reg.scala 15:16]
  reg [7:0] r_24_1; // @[Reg.scala 15:16]
  reg [7:0] r_25_0; // @[Reg.scala 15:16]
  reg [7:0] r_25_1; // @[Reg.scala 15:16]
  reg  r_26_0; // @[Reg.scala 15:16]
  reg  r_27_0; // @[Reg.scala 15:16]
  reg  r_28_0; // @[Reg.scala 15:16]
  reg  r_29_0; // @[Reg.scala 15:16]
  wire [1:0] _T_141 = ~io_req_bits_pe_control_dataflow ? 2'h3 : 2'h2; // @[MeshWithDelays.scala 218:55]
  wire [2:0] _GEN_88 = {{1'd0}, _T_141}; // @[Util.scala 13:22]
  wire [2:0] _T_147 = 3'h4 - _GEN_88; // @[Util.scala 13:22]
  wire [2:0] _T_149 = _T_147 + 3'h1; // @[Util.scala 13:26]
  wire [2:0] _T_156 = _GEN_88 - _T_24; // @[Util.scala 13:48]
  wire [2:0] _T_158 = _T_156 - 3'h1; // @[Util.scala 13:62]
  wire [2:0] _T_160 = matmul_id + _GEN_88; // @[Util.scala 13:71]
  wire  _T_181 = io_req_bits_flush == 2'h0; // @[MeshWithDelays.scala 222:57]
  reg [2:0] r_30_0; // @[Reg.scala 15:16]
  reg [2:0] r_31_0; // @[Reg.scala 15:16]
  wire [2:0] out_matmul_id = r_31_0;
  wire  _T_183 = out_matmul_id == tagq_io_deq_bits_id; // @[MeshWithDelays.scala 232:62]
  wire  _T_186 = io_resp_valid & io_resp_bits_last; // @[MeshWithDelays.scala 236:38]
  wire  _T_192 = out_matmul_id == total_rows_q_io_deq_bits_id; // @[MeshWithDelays.scala 244:77]
  AlwaysOutTransposer transposer ( // @[MeshWithDelays.scala 154:26]
    .clock(transposer_clock),
    .reset(transposer_reset),
    .io_inRow_ready(transposer_io_inRow_ready),
    .io_inRow_valid(transposer_io_inRow_valid),
    .io_inRow_bits_0(transposer_io_inRow_bits_0),
    .io_inRow_bits_1(transposer_io_inRow_bits_1),
    .io_inRow_bits_2(transposer_io_inRow_bits_2),
    .io_inRow_bits_3(transposer_io_inRow_bits_3),
    .io_outCol_bits_0(transposer_io_outCol_bits_0),
    .io_outCol_bits_1(transposer_io_outCol_bits_1),
    .io_outCol_bits_2(transposer_io_outCol_bits_2),
    .io_outCol_bits_3(transposer_io_outCol_bits_3)
  );
  Mesh mesh ( // @[MeshWithDelays.scala 166:20]
    .clock(mesh_clock),
    .io_in_a_0_0(mesh_io_in_a_0_0),
    .io_in_a_0_1(mesh_io_in_a_0_1),
    .io_in_a_1_0(mesh_io_in_a_1_0),
    .io_in_a_1_1(mesh_io_in_a_1_1),
    .io_in_b_0_0(mesh_io_in_b_0_0),
    .io_in_b_0_1(mesh_io_in_b_0_1),
    .io_in_b_1_0(mesh_io_in_b_1_0),
    .io_in_b_1_1(mesh_io_in_b_1_1),
    .io_in_d_0_0(mesh_io_in_d_0_0),
    .io_in_d_0_1(mesh_io_in_d_0_1),
    .io_in_d_1_0(mesh_io_in_d_1_0),
    .io_in_d_1_1(mesh_io_in_d_1_1),
    .io_in_control_0_0_dataflow(mesh_io_in_control_0_0_dataflow),
    .io_in_control_0_0_propagate(mesh_io_in_control_0_0_propagate),
    .io_in_control_0_0_shift(mesh_io_in_control_0_0_shift),
    .io_in_control_0_1_dataflow(mesh_io_in_control_0_1_dataflow),
    .io_in_control_0_1_propagate(mesh_io_in_control_0_1_propagate),
    .io_in_control_0_1_shift(mesh_io_in_control_0_1_shift),
    .io_in_control_1_0_dataflow(mesh_io_in_control_1_0_dataflow),
    .io_in_control_1_0_propagate(mesh_io_in_control_1_0_propagate),
    .io_in_control_1_0_shift(mesh_io_in_control_1_0_shift),
    .io_in_control_1_1_dataflow(mesh_io_in_control_1_1_dataflow),
    .io_in_control_1_1_propagate(mesh_io_in_control_1_1_propagate),
    .io_in_control_1_1_shift(mesh_io_in_control_1_1_shift),
    .io_in_id_0_0(mesh_io_in_id_0_0),
    .io_in_id_0_1(mesh_io_in_id_0_1),
    .io_in_id_1_0(mesh_io_in_id_1_0),
    .io_in_id_1_1(mesh_io_in_id_1_1),
    .io_in_last_0_0(mesh_io_in_last_0_0),
    .io_in_last_0_1(mesh_io_in_last_0_1),
    .io_in_last_1_0(mesh_io_in_last_1_0),
    .io_in_last_1_1(mesh_io_in_last_1_1),
    .io_out_b_0_0(mesh_io_out_b_0_0),
    .io_out_b_0_1(mesh_io_out_b_0_1),
    .io_out_b_1_0(mesh_io_out_b_1_0),
    .io_out_b_1_1(mesh_io_out_b_1_1),
    .io_out_c_0_0(mesh_io_out_c_0_0),
    .io_out_c_0_1(mesh_io_out_c_0_1),
    .io_out_c_1_0(mesh_io_out_c_1_0),
    .io_out_c_1_1(mesh_io_out_c_1_1),
    .io_in_valid_0_0(mesh_io_in_valid_0_0),
    .io_in_valid_0_1(mesh_io_in_valid_0_1),
    .io_in_valid_1_0(mesh_io_in_valid_1_0),
    .io_in_valid_1_1(mesh_io_in_valid_1_1),
    .io_out_valid_0_0(mesh_io_out_valid_0_0),
    .io_out_control_0_0_dataflow(mesh_io_out_control_0_0_dataflow),
    .io_out_id_0_0(mesh_io_out_id_0_0),
    .io_out_last_0_0(mesh_io_out_last_0_0)
  );
  TagQueue tagq ( // @[MeshWithDelays.scala 221:20]
    .clock(tagq_clock),
    .reset(tagq_reset),
    .io_enq_ready(tagq_io_enq_ready),
    .io_enq_valid(tagq_io_enq_valid),
    .io_enq_bits_tag(tagq_io_enq_bits_tag),
    .io_enq_bits_id(tagq_io_enq_bits_id),
    .io_deq_ready(tagq_io_deq_ready),
    .io_deq_valid(tagq_io_deq_valid),
    .io_deq_bits_tag(tagq_io_deq_bits_tag),
    .io_deq_bits_id(tagq_io_deq_bits_id),
    .io_all_0_tag(tagq_io_all_0_tag),
    .io_all_1_tag(tagq_io_all_1_tag),
    .io_all_2_tag(tagq_io_all_2_tag),
    .io_all_3_tag(tagq_io_all_3_tag),
    .io_all_4_tag(tagq_io_all_4_tag),
    .io_all_5_tag(tagq_io_all_5_tag)
  );
  Queue total_rows_q ( // @[MeshWithDelays.scala 238:28]
    .clock(total_rows_q_clock),
    .reset(total_rows_q_reset),
    .io_enq_ready(total_rows_q_io_enq_ready),
    .io_enq_valid(total_rows_q_io_enq_valid),
    .io_enq_bits_id(total_rows_q_io_enq_bits_id),
    .io_enq_bits_total_rows(total_rows_q_io_enq_bits_total_rows),
    .io_deq_ready(total_rows_q_io_deq_ready),
    .io_deq_valid(total_rows_q_io_deq_valid),
    .io_deq_bits_id(total_rows_q_io_deq_bits_id),
    .io_deq_bits_total_rows(total_rows_q_io_deq_bits_total_rows)
  );
  assign io_a_ready = ~a_written | input_next_row_into_spatial_array | io_req_ready; // @[MeshWithDelays.scala 142:65]
  assign io_b_ready = ~b_written | input_next_row_into_spatial_array | io_req_ready; // @[MeshWithDelays.scala 143:65]
  assign io_d_ready = ~d_written | input_next_row_into_spatial_array | io_req_ready; // @[MeshWithDelays.scala 144:65]
  assign io_req_ready = (_T_80 | last_fire) & tagq_io_enq_ready & total_rows_q_io_enq_ready; // @[MeshWithDelays.scala 249:66]
  assign io_resp_valid = r_27_0; // @[MeshWithDelays.scala 200:17]
  assign io_resp_bits_data_0_0 = r_25_0; // @[MeshWithDelays.scala 198:21]
  assign io_resp_bits_data_0_1 = r_25_1; // @[MeshWithDelays.scala 198:21]
  assign io_resp_bits_data_1_0 = ~mesh_io_out_control_0_0_dataflow ? $signed(mesh_io_out_c_1_0) : $signed(
    mesh_io_out_b_1_0); // @[MeshWithDelays.scala 198:35]
  assign io_resp_bits_data_1_1 = ~mesh_io_out_control_0_0_dataflow ? $signed(mesh_io_out_c_1_1) : $signed(
    mesh_io_out_b_1_1); // @[MeshWithDelays.scala 198:35]
  assign io_resp_bits_total_rows = total_rows_q_io_deq_valid & out_matmul_id == total_rows_q_io_deq_bits_id ?
    total_rows_q_io_deq_bits_total_rows : 3'h4; // @[MeshWithDelays.scala 244:33]
  assign io_resp_bits_tag = tagq_io_deq_valid & out_matmul_id == tagq_io_deq_bits_id ? tagq_io_deq_bits_tag : 32'h0; // @[MeshWithDelays.scala 232:26]
  assign io_resp_bits_last = r_29_0; // @[MeshWithDelays.scala 203:21]
  assign io_tags_in_progress_0 = tagq_io_all_0_tag; // @[MeshWithDelays.scala 250:23]
  assign io_tags_in_progress_1 = tagq_io_all_1_tag; // @[MeshWithDelays.scala 250:23]
  assign io_tags_in_progress_2 = tagq_io_all_2_tag; // @[MeshWithDelays.scala 250:23]
  assign io_tags_in_progress_3 = tagq_io_all_3_tag; // @[MeshWithDelays.scala 250:23]
  assign io_tags_in_progress_4 = tagq_io_all_4_tag; // @[MeshWithDelays.scala 250:23]
  assign io_tags_in_progress_5 = tagq_io_all_5_tag; // @[MeshWithDelays.scala 250:23]
  assign transposer_clock = clock;
  assign transposer_reset = reset;
  assign transposer_io_inRow_valid = ~pause & (a_is_from_transposer | b_is_from_transposer | d_is_from_transposer); // @[MeshWithDelays.scala 156:39]
  assign transposer_io_inRow_bits_0 = b_is_from_transposer ? $signed(b_buf_0_0) : $signed(_T_90_0); // @[Mux.scala 98:16]
  assign transposer_io_inRow_bits_1 = b_is_from_transposer ? $signed(b_buf_0_1) : $signed(_T_90_1); // @[Mux.scala 98:16]
  assign transposer_io_inRow_bits_2 = b_is_from_transposer ? $signed(b_buf_1_0) : $signed(_T_90_2); // @[Mux.scala 98:16]
  assign transposer_io_inRow_bits_3 = b_is_from_transposer ? $signed(b_buf_1_1) : $signed(_T_90_3); // @[Mux.scala 98:16]
  assign mesh_clock = clock;
  assign mesh_io_in_a_0_0 = a_is_from_transposer ? $signed(_T_98) : $signed(a_buf_0_0); // @[MeshWithDelays.scala 169:34]
  assign mesh_io_in_a_0_1 = a_is_from_transposer ? $signed(_T_100) : $signed(a_buf_0_1); // @[MeshWithDelays.scala 169:34]
  assign mesh_io_in_a_1_0 = r_1_0; // @[MeshWithDelays.scala 174:16]
  assign mesh_io_in_a_1_1 = r_1_1; // @[MeshWithDelays.scala 174:16]
  assign mesh_io_in_b_0_0 = b_is_from_transposer ? $signed(_T_98) : $signed(b_buf_0_0); // @[MeshWithDelays.scala 170:34]
  assign mesh_io_in_b_0_1 = b_is_from_transposer ? $signed(_T_100) : $signed(b_buf_0_1); // @[MeshWithDelays.scala 170:34]
  assign mesh_io_in_b_1_0 = r_3_0; // @[MeshWithDelays.scala 175:16]
  assign mesh_io_in_b_1_1 = r_3_1; // @[MeshWithDelays.scala 175:16]
  assign mesh_io_in_d_0_0 = d_is_from_transposer ? $signed(_T_126) : $signed(d_buf_0_0); // @[MeshWithDelays.scala 171:34]
  assign mesh_io_in_d_0_1 = d_is_from_transposer ? $signed(_T_128) : $signed(d_buf_0_1); // @[MeshWithDelays.scala 171:34]
  assign mesh_io_in_d_1_0 = r_5_0; // @[MeshWithDelays.scala 176:16]
  assign mesh_io_in_d_1_1 = r_5_1; // @[MeshWithDelays.scala 176:16]
  assign mesh_io_in_control_0_0_dataflow = req_bits_pe_control_dataflow; // @[MeshWithDelays.scala 179:27]
  assign mesh_io_in_control_0_0_propagate = in_prop; // @[MeshWithDelays.scala 180:28]
  assign mesh_io_in_control_0_0_shift = result_shift; // @[MeshWithDelays.scala 184:26]
  assign mesh_io_in_control_0_1_dataflow = req_bits_pe_control_dataflow; // @[MeshWithDelays.scala 179:27]
  assign mesh_io_in_control_0_1_propagate = in_prop; // @[MeshWithDelays.scala 180:28]
  assign mesh_io_in_control_0_1_shift = result_shift; // @[MeshWithDelays.scala 184:26]
  assign mesh_io_in_control_1_0_dataflow = r_7; // @[MeshWithDelays.scala 179:27]
  assign mesh_io_in_control_1_0_propagate = r_11; // @[MeshWithDelays.scala 180:28]
  assign mesh_io_in_control_1_0_shift = r_15; // @[MeshWithDelays.scala 184:26]
  assign mesh_io_in_control_1_1_dataflow = r_9; // @[MeshWithDelays.scala 179:27]
  assign mesh_io_in_control_1_1_propagate = r_13; // @[MeshWithDelays.scala 180:28]
  assign mesh_io_in_control_1_1_shift = r_17; // @[MeshWithDelays.scala 184:26]
  assign mesh_io_in_id_0_0 = matmul_id; // @[MeshWithDelays.scala 190:60 MeshWithDelays.scala 190:60]
  assign mesh_io_in_id_0_1 = matmul_id; // @[MeshWithDelays.scala 190:60 MeshWithDelays.scala 190:60]
  assign mesh_io_in_id_1_0 = r_21_0; // @[MeshWithDelays.scala 191:17]
  assign mesh_io_in_id_1_1 = r_21_1; // @[MeshWithDelays.scala 191:17]
  assign mesh_io_in_last_0_0 = _GEN_85 == _T_8 & input_next_row_into_spatial_array; // @[MeshWithDelays.scala 111:54]
  assign mesh_io_in_last_0_1 = _GEN_85 == _T_8 & input_next_row_into_spatial_array; // @[MeshWithDelays.scala 111:54]
  assign mesh_io_in_last_1_0 = r_23_0; // @[MeshWithDelays.scala 194:19]
  assign mesh_io_in_last_1_1 = r_23_1; // @[MeshWithDelays.scala 194:19]
  assign mesh_io_in_valid_0_0 = ~pause; // @[MeshWithDelays.scala 187:84]
  assign mesh_io_in_valid_0_1 = ~pause; // @[MeshWithDelays.scala 187:84]
  assign mesh_io_in_valid_1_0 = r_19_0; // @[MeshWithDelays.scala 188:20]
  assign mesh_io_in_valid_1_1 = r_19_1; // @[MeshWithDelays.scala 188:20]
  assign tagq_clock = clock;
  assign tagq_reset = reset;
  assign tagq_io_enq_valid = _T_10 & io_req_bits_flush == 2'h0; // @[MeshWithDelays.scala 222:36]
  assign tagq_io_enq_bits_tag = io_req_bits_tag; // @[MeshWithDelays.scala 223:24]
  assign tagq_io_enq_bits_id = matmul_id >= _T_149 & _T_141 != 2'h0 ? _T_158 : _T_160; // @[Util.scala 13:10]
  assign tagq_io_deq_ready = io_resp_valid & io_resp_bits_last & _T_183; // @[MeshWithDelays.scala 236:59]
  assign total_rows_q_clock = clock;
  assign total_rows_q_reset = reset;
  assign total_rows_q_io_enq_valid = _T_10 & _T_181; // @[MeshWithDelays.scala 239:44]
  assign total_rows_q_io_enq_bits_id = matmul_id >= _T_19 ? _T_28 : _T_30; // @[Util.scala 13:10]
  assign total_rows_q_io_enq_bits_total_rows = io_req_bits_total_rows; // @[MeshWithDelays.scala 241:39]
  assign total_rows_q_io_deq_ready = _T_186 & _T_192; // @[MeshWithDelays.scala 247:67]
  always @(posedge clock) begin
    if (reset) begin // @[MeshWithDelays.scala 252:25]
      req_valid <= 1'h0; // @[MeshWithDelays.scala 253:15]
    end else begin
      req_valid <= _GEN_14;
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      req_bits_pe_control_dataflow <= io_req_bits_pe_control_dataflow; // @[Util.scala 135:12]
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      req_bits_pe_control_shift <= io_req_bits_pe_control_shift; // @[Util.scala 135:12]
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      req_bits_a_transpose <= io_req_bits_a_transpose; // @[Util.scala 135:12]
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      req_bits_bd_transpose <= io_req_bits_bd_transpose; // @[Util.scala 135:12]
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      req_bits_total_rows <= io_req_bits_total_rows; // @[Util.scala 135:12]
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      req_bits_flush <= io_req_bits_flush; // @[Util.scala 135:12]
    end else if (last_fire) begin // @[MeshWithDelays.scala 117:26]
      req_bits_flush <= _T_34; // @[MeshWithDelays.scala 119:20]
    end
    if (reset) begin // @[MeshWithDelays.scala 94:26]
      matmul_id <= 3'h0; // @[MeshWithDelays.scala 94:26]
    end else if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      if (matmul_id >= _T_19) begin // @[Util.scala 13:10]
        matmul_id <= _T_28;
      end else begin
        matmul_id <= _T_30;
      end
    end
    if (reset) begin // @[MeshWithDelays.scala 97:29]
      fire_counter <= 2'h0; // @[MeshWithDelays.scala 97:29]
    end else begin
      fire_counter <= _GEN_28[1:0];
    end
    if (_T) begin // @[Reg.scala 16:19]
      a_buf_0_0 <= io_a_bits_0_0; // @[Reg.scala 16:23]
    end
    if (_T) begin // @[Reg.scala 16:19]
      a_buf_0_1 <= io_a_bits_0_1; // @[Reg.scala 16:23]
    end
    if (_T) begin // @[Reg.scala 16:19]
      a_buf_1_0 <= io_a_bits_1_0; // @[Reg.scala 16:23]
    end
    if (_T) begin // @[Reg.scala 16:19]
      a_buf_1_1 <= io_a_bits_1_1; // @[Reg.scala 16:23]
    end
    if (_T_1) begin // @[Reg.scala 16:19]
      b_buf_0_0 <= io_b_bits_0_0; // @[Reg.scala 16:23]
    end
    if (_T_1) begin // @[Reg.scala 16:19]
      b_buf_0_1 <= io_b_bits_0_1; // @[Reg.scala 16:23]
    end
    if (_T_1) begin // @[Reg.scala 16:19]
      b_buf_1_0 <= io_b_bits_1_0; // @[Reg.scala 16:23]
    end
    if (_T_1) begin // @[Reg.scala 16:19]
      b_buf_1_1 <= io_b_bits_1_1; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      d_buf_0_0 <= io_d_bits_0_0; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      d_buf_0_1 <= io_d_bits_0_1; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      d_buf_1_0 <= io_d_bits_1_0; // @[Reg.scala 16:23]
    end
    if (_T_2) begin // @[Reg.scala 16:19]
      d_buf_1_1 <= io_d_bits_1_1; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[MeshWithDelays.scala 103:26]
      a_written <= 1'h0; // @[MeshWithDelays.scala 103:26]
    end else begin
      a_written <= _GEN_29;
    end
    if (reset) begin // @[MeshWithDelays.scala 104:26]
      b_written <= 1'h0; // @[MeshWithDelays.scala 104:26]
    end else begin
      b_written <= _GEN_30;
    end
    if (reset) begin // @[MeshWithDelays.scala 105:26]
      d_written <= 1'h0; // @[MeshWithDelays.scala 105:26]
    end else begin
      d_written <= _GEN_31;
    end
    if (_T_10) begin // @[MeshWithDelays.scala 113:22]
      in_prop <= io_req_bits_pe_control_propagate ^ in_prop; // @[MeshWithDelays.scala 115:13]
    end
    if (a_is_from_transposer) begin // @[MeshWithDelays.scala 169:34]
      r__0 <= _T_102;
    end else begin
      r__0 <= a_buf_1_0;
    end
    if (a_is_from_transposer) begin // @[MeshWithDelays.scala 169:34]
      r__1 <= _T_104;
    end else begin
      r__1 <= a_buf_1_1;
    end
    r_1_0 <= r__0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_1_1 <= r__1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    if (b_is_from_transposer) begin // @[MeshWithDelays.scala 170:34]
      r_2_0 <= _T_102;
    end else begin
      r_2_0 <= b_buf_1_0;
    end
    if (b_is_from_transposer) begin // @[MeshWithDelays.scala 170:34]
      r_2_1 <= _T_104;
    end else begin
      r_2_1 <= b_buf_1_1;
    end
    r_3_0 <= r_2_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_3_1 <= r_2_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    if (d_is_from_transposer) begin // @[MeshWithDelays.scala 171:34]
      r_4_0 <= _T_130;
    end else begin
      r_4_0 <= d_buf_1_0;
    end
    if (d_is_from_transposer) begin // @[MeshWithDelays.scala 171:34]
      r_4_1 <= _T_132;
    end else begin
      r_4_1 <= d_buf_1_1;
    end
    r_5_0 <= r_4_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_5_1 <= r_4_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_6 <= req_bits_pe_control_dataflow; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_7 <= r_6; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_8 <= req_bits_pe_control_dataflow; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_9 <= r_8; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_10 <= in_prop; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_11 <= r_10; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_12 <= in_prop; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_13 <= r_12; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    result_shift <= req_bits_pe_control_shift; // @[MeshWithDelays.scala 182:29]
    r_14 <= result_shift; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_15 <= r_14; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_16 <= result_shift; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_17 <= r_16; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_18_0 <= ~pause; // @[MeshWithDelays.scala 187:84]
    r_18_1 <= ~pause; // @[MeshWithDelays.scala 187:84]
    r_19_0 <= r_18_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_19_1 <= r_18_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_20_0 <= matmul_id; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_20_1 <= matmul_id; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_21_0 <= r_20_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_21_1 <= r_20_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_22_0 <= _GEN_85 == _T_8 & input_next_row_into_spatial_array; // @[MeshWithDelays.scala 111:54]
    r_22_1 <= _GEN_85 == _T_8 & input_next_row_into_spatial_array; // @[MeshWithDelays.scala 111:54]
    r_23_0 <= r_22_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_23_1 <= r_22_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    if (~mesh_io_out_control_0_0_dataflow) begin // @[MeshWithDelays.scala 198:35]
      r_24_0 <= mesh_io_out_c_0_0;
    end else begin
      r_24_0 <= mesh_io_out_b_0_0;
    end
    if (~mesh_io_out_control_0_0_dataflow) begin // @[MeshWithDelays.scala 198:35]
      r_24_1 <= mesh_io_out_c_0_1;
    end else begin
      r_24_1 <= mesh_io_out_b_0_1;
    end
    r_25_0 <= r_24_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_25_1 <= r_24_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_26_0 <= mesh_io_out_valid_0_0; // @[MeshWithDelays.scala 78:26 MeshWithDelays.scala 78:26]
    r_27_0 <= r_26_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_28_0 <= mesh_io_out_last_0_0; // @[MeshWithDelays.scala 78:26 MeshWithDelays.scala 78:26]
    r_29_0 <= r_28_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_30_0 <= mesh_io_out_id_0_0; // @[MeshWithDelays.scala 78:26 MeshWithDelays.scala 78:26]
    r_31_0 <= r_30_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (input_next_row_into_spatial_array & ~(3'h1 <= _T_8 | _T_8 == 3'h0 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: cannot wrapAdd when n is larger than max, unless max is 0\n    at Util.scala:19 assert(n <= max || max === 0.U, \"cannot wrapAdd when n is larger than max, unless max is 0\")\n"
            ); // @[Util.scala 19:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (input_next_row_into_spatial_array & ~(3'h1 <= _T_8 | _T_8 == 3'h0 | reset)) begin
          $fatal; // @[Util.scala 19:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(req_valid | ~input_next_row_into_spatial_array | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at MeshWithDelays.scala:146 assert(req.valid || !input_next_row_into_spatial_array)\n"
            ); // @[MeshWithDelays.scala 146:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(req_valid | ~input_next_row_into_spatial_array | reset)) begin
          $fatal; // @[MeshWithDelays.scala 146:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(_T_10 & ~tagq_io_enq_ready & _T_181) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at MeshWithDelays.scala:256 assert(!(io.req.fire && !tagq.io.enq.ready && io.req.bits.flush === 0.U))\n"
            ); // @[MeshWithDelays.scala 256:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(_T_10 & ~tagq_io_enq_ready & _T_181) | reset)) begin
          $fatal; // @[MeshWithDelays.scala 256:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  req_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  req_bits_pe_control_dataflow = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  req_bits_pe_control_shift = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  req_bits_a_transpose = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  req_bits_bd_transpose = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  req_bits_total_rows = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  req_bits_flush = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  matmul_id = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  fire_counter = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  a_buf_0_0 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  a_buf_0_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  a_buf_1_0 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  a_buf_1_1 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  b_buf_0_0 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  b_buf_0_1 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  b_buf_1_0 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  b_buf_1_1 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  d_buf_0_0 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  d_buf_0_1 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  d_buf_1_0 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  d_buf_1_1 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  a_written = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  b_written = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  d_written = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  in_prop = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r__0 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  r__1 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  r_1_0 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  r_1_1 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  r_2_0 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  r_2_1 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  r_3_0 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  r_3_1 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  r_4_0 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  r_4_1 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  r_5_0 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  r_5_1 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  r_6 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_7 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_8 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_9 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_10 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_11 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_12 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_13 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  result_shift = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  r_14 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  r_15 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  r_16 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  r_17 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  r_18_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  r_18_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_19_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_19_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r_20_0 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  r_20_1 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  r_21_0 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  r_21_1 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  r_22_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_22_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  r_23_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_23_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_24_0 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  r_24_1 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  r_25_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  r_25_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  r_26_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r_27_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  r_28_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  r_29_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  r_30_0 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  r_31_0 = _RAND_71[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
